module sha256_unrolled_pipelined (clk,
    ready,
    reset,
    hashvalue,
    message);
 input clk;
 output ready;
 input reset;
 output [255:0] hashvalue;
 input [0:511] message;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire net629;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire net1;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire net551;
 wire net550;
 wire net549;
 wire net548;
 wire net547;
 wire net546;
 wire net545;
 wire net544;
 wire net543;
 wire _02714_;
 wire net542;
 wire net541;
 wire _02717_;
 wire _02718_;
 wire net540;
 wire net539;
 wire net538;
 wire _02722_;
 wire net537;
 wire net536;
 wire net535;
 wire net534;
 wire net533;
 wire _02728_;
 wire _02729_;
 wire net532;
 wire net531;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire net530;
 wire net529;
 wire _02738_;
 wire net528;
 wire net527;
 wire net526;
 wire _02742_;
 wire net525;
 wire net524;
 wire _02745_;
 wire net523;
 wire net522;
 wire _02748_;
 wire net521;
 wire net520;
 wire _02751_;
 wire net519;
 wire net518;
 wire _02754_;
 wire net517;
 wire _02756_;
 wire net516;
 wire net515;
 wire _02759_;
 wire net514;
 wire net513;
 wire _02762_;
 wire net512;
 wire net511;
 wire _02765_;
 wire net510;
 wire net509;
 wire _02768_;
 wire net508;
 wire _02770_;
 wire net507;
 wire _02772_;
 wire net506;
 wire net505;
 wire _02775_;
 wire _02776_;
 wire net504;
 wire net503;
 wire _02779_;
 wire net502;
 wire net501;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire net500;
 wire net499;
 wire net498;
 wire net497;
 wire net496;
 wire net495;
 wire net494;
 wire net493;
 wire net492;
 wire _02799_;
 wire net491;
 wire net490;
 wire net489;
 wire net488;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire net487;
 wire net486;
 wire net485;
 wire net484;
 wire net483;
 wire _02812_;
 wire _02813_;
 wire net482;
 wire net481;
 wire net480;
 wire net479;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire net478;
 wire net477;
 wire _02824_;
 wire net476;
 wire net475;
 wire _02827_;
 wire net474;
 wire net473;
 wire _02830_;
 wire net472;
 wire net471;
 wire _02833_;
 wire net470;
 wire net469;
 wire _02836_;
 wire net468;
 wire net467;
 wire _02839_;
 wire _02840_;
 wire net466;
 wire _02842_;
 wire net465;
 wire net464;
 wire _02845_;
 wire net463;
 wire net462;
 wire _02848_;
 wire net461;
 wire net460;
 wire _02851_;
 wire net459;
 wire _02853_;
 wire net458;
 wire net457;
 wire _02856_;
 wire net456;
 wire net455;
 wire _02859_;
 wire net454;
 wire _02861_;
 wire net453;
 wire _02863_;
 wire net452;
 wire net451;
 wire _02866_;
 wire net450;
 wire net449;
 wire _02869_;
 wire net448;
 wire net447;
 wire _02872_;
 wire net446;
 wire net445;
 wire _02875_;
 wire net444;
 wire net443;
 wire _02878_;
 wire net442;
 wire net441;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire net440;
 wire net439;
 wire net438;
 wire net437;
 wire net436;
 wire net435;
 wire net434;
 wire net433;
 wire _02892_;
 wire net432;
 wire net431;
 wire net430;
 wire net429;
 wire _02897_;
 wire net428;
 wire net427;
 wire _02900_;
 wire net426;
 wire net425;
 wire net424;
 wire _02904_;
 wire net423;
 wire net422;
 wire net421;
 wire net420;
 wire net419;
 wire _02910_;
 wire net418;
 wire net417;
 wire _02913_;
 wire net416;
 wire net415;
 wire _02916_;
 wire net414;
 wire net413;
 wire _02919_;
 wire net412;
 wire net411;
 wire _02922_;
 wire net410;
 wire net409;
 wire _02925_;
 wire net408;
 wire net407;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire net406;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire net405;
 wire _02947_;
 wire _02948_;
 wire net404;
 wire _02950_;
 wire net403;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire net402;
 wire net401;
 wire _02980_;
 wire _02981_;
 wire net400;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire net399;
 wire net398;
 wire _02989_;
 wire net397;
 wire net396;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire net395;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire net394;
 wire net393;
 wire net392;
 wire net391;
 wire net390;
 wire net389;
 wire net388;
 wire net387;
 wire _03026_;
 wire net386;
 wire net385;
 wire net384;
 wire net383;
 wire _03031_;
 wire net382;
 wire net381;
 wire _03034_;
 wire net380;
 wire net379;
 wire net378;
 wire _03038_;
 wire net377;
 wire net376;
 wire net375;
 wire net374;
 wire net373;
 wire _03044_;
 wire net372;
 wire net371;
 wire _03047_;
 wire net370;
 wire net369;
 wire _03050_;
 wire net368;
 wire net367;
 wire _03053_;
 wire net366;
 wire net365;
 wire _03056_;
 wire net364;
 wire net363;
 wire _03059_;
 wire net362;
 wire net361;
 wire net360;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire net359;
 wire _03072_;
 wire net358;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire net357;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire net356;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire net355;
 wire net354;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire net353;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire net352;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire net351;
 wire net350;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire net349;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire net348;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire net347;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire net346;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire net345;
 wire _03283_;
 wire _03284_;
 wire net344;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire net343;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire net342;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire net341;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire net340;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire net339;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire net338;
 wire _03425_;
 wire net337;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire net336;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire net335;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire net334;
 wire _03484_;
 wire net333;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire net332;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire net331;
 wire _03537_;
 wire net330;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire net329;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire net328;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire net327;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire net326;
 wire _03604_;
 wire net325;
 wire _03606_;
 wire net324;
 wire _03608_;
 wire net323;
 wire _03610_;
 wire net322;
 wire _03612_;
 wire net321;
 wire _03614_;
 wire net320;
 wire _03616_;
 wire net319;
 wire _03618_;
 wire net318;
 wire _03620_;
 wire net317;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire net316;
 wire net315;
 wire _03670_;
 wire net314;
 wire _03672_;
 wire net313;
 wire _03674_;
 wire net312;
 wire _03676_;
 wire _03677_;
 wire net311;
 wire _03679_;
 wire net310;
 wire _03681_;
 wire net309;
 wire _03683_;
 wire net308;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire net307;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire net306;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire net305;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire net304;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire net303;
 wire net302;
 wire _03781_;
 wire net301;
 wire net300;
 wire _03784_;
 wire net299;
 wire net298;
 wire _03787_;
 wire net297;
 wire net296;
 wire _03790_;
 wire net295;
 wire net294;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire net293;
 wire net292;
 wire _03798_;
 wire net291;
 wire net290;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire net289;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire net288;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire net287;
 wire _03853_;
 wire net286;
 wire net285;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03872_;
 wire _03873_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire net1141;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire net1140;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire net1139;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire net1138;
 wire _03968_;
 wire net1137;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire net1136;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire net1135;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire net1134;
 wire _04005_;
 wire net1133;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire net1129;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire net1128;
 wire _04036_;
 wire net1127;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire net1125;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire net1124;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire net1123;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire net1122;
 wire _04081_;
 wire net1121;
 wire _04083_;
 wire net1120;
 wire _04085_;
 wire net1119;
 wire _04087_;
 wire net1118;
 wire _04089_;
 wire net1117;
 wire _04091_;
 wire net1116;
 wire _04093_;
 wire net1115;
 wire _04095_;
 wire net1110;
 wire _04097_;
 wire net1105;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire net1104;
 wire net1103;
 wire _04125_;
 wire net1102;
 wire _04127_;
 wire net1101;
 wire _04129_;
 wire net1098;
 wire _04131_;
 wire _04132_;
 wire net1097;
 wire _04134_;
 wire net1096;
 wire _04136_;
 wire net1095;
 wire _04138_;
 wire net1094;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire net1093;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire net1114;
 wire net1113;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire net1112;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire net1111;
 wire net1108;
 wire net1107;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire net1100;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire net1099;
 wire _04389_;
 wire net1092;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire net1091;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire net1090;
 wire _04439_;
 wire net1089;
 wire net1088;
 wire _04442_;
 wire net1087;
 wire net1086;
 wire net1085;
 wire _04446_;
 wire net1084;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire net1083;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire net1082;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire net1081;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire net1080;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire net1079;
 wire net1078;
 wire net1077;
 wire net1076;
 wire net1075;
 wire _04784_;
 wire net1074;
 wire _04786_;
 wire net1073;
 wire net1072;
 wire net1071;
 wire _04790_;
 wire net1070;
 wire net1069;
 wire _04793_;
 wire _04794_;
 wire net1068;
 wire _04796_;
 wire _04797_;
 wire net1067;
 wire net1066;
 wire _04800_;
 wire _04801_;
 wire net1065;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire net1064;
 wire _04807_;
 wire _04808_;
 wire net1063;
 wire _04810_;
 wire net1062;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire net1061;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire net1060;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire net1059;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire net1058;
 wire _04845_;
 wire net1057;
 wire net1056;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire net1055;
 wire _04854_;
 wire net1054;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire net1053;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire net1052;
 wire net1051;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire net1050;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire net1049;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire net1048;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire net1047;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire net1046;
 wire _04913_;
 wire net1045;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire net1044;
 wire _04925_;
 wire net1043;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire net1042;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire net1041;
 wire _04941_;
 wire net1040;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire clknet_5_31__leaf_clk;
 wire _04953_;
 wire clknet_5_30__leaf_clk;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire _04963_;
 wire clknet_5_27__leaf_clk;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire clknet_5_26__leaf_clk;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire clknet_5_25__leaf_clk;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire clknet_5_24__leaf_clk;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire clknet_5_23__leaf_clk;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire clknet_5_22__leaf_clk;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire clknet_5_21__leaf_clk;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire clknet_5_20__leaf_clk;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire clknet_5_19__leaf_clk;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire clknet_5_18__leaf_clk;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire clknet_5_17__leaf_clk;
 wire _05062_;
 wire _05063_;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire clknet_5_12__leaf_clk;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire clknet_5_11__leaf_clk;
 wire _05080_;
 wire _05081_;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire clknet_5_6__leaf_clk;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire clknet_5_5__leaf_clk;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire clknet_5_4__leaf_clk;
 wire _05118_;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire _05121_;
 wire _05122_;
 wire clknet_5_1__leaf_clk;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire clknet_5_0__leaf_clk;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire clknet_2_3_0_clk;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire clknet_2_2_0_clk;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire clknet_2_1_0_clk;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire clknet_2_0_0_clk;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire clknet_0_clk;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire clknet_leaf_290_clk;
 wire _05175_;
 wire clknet_leaf_289_clk;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire clknet_leaf_288_clk;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire clknet_leaf_287_clk;
 wire clknet_leaf_286_clk;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire clknet_leaf_285_clk;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire clknet_leaf_284_clk;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire clknet_leaf_283_clk;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire clknet_leaf_282_clk;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire clknet_leaf_281_clk;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire clknet_leaf_280_clk;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire clknet_leaf_279_clk;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire clknet_leaf_278_clk;
 wire _05269_;
 wire clknet_leaf_277_clk;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire clknet_leaf_276_clk;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire clknet_leaf_275_clk;
 wire clknet_leaf_274_clk;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire clknet_leaf_273_clk;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire clknet_leaf_272_clk;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire clknet_leaf_271_clk;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire clknet_leaf_270_clk;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire clknet_leaf_269_clk;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire clknet_leaf_268_clk;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire clknet_leaf_267_clk;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire clknet_leaf_266_clk;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire clknet_leaf_265_clk;
 wire _05382_;
 wire clknet_leaf_264_clk;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire clknet_leaf_263_clk;
 wire _05432_;
 wire _05433_;
 wire clknet_leaf_262_clk;
 wire _05435_;
 wire clknet_leaf_261_clk;
 wire clknet_leaf_260_clk;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire clknet_leaf_259_clk;
 wire _05447_;
 wire _05448_;
 wire clknet_leaf_258_clk;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire clknet_leaf_257_clk;
 wire _05459_;
 wire _05460_;
 wire clknet_leaf_256_clk;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire clknet_leaf_255_clk;
 wire clknet_leaf_254_clk;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire clknet_leaf_253_clk;
 wire _05488_;
 wire clknet_leaf_252_clk;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire clknet_leaf_251_clk;
 wire _05500_;
 wire clknet_leaf_250_clk;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire clknet_leaf_249_clk;
 wire clknet_leaf_248_clk;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire clknet_leaf_247_clk;
 wire _05518_;
 wire clknet_leaf_246_clk;
 wire clknet_leaf_245_clk;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire clknet_leaf_244_clk;
 wire _05530_;
 wire _05531_;
 wire clknet_leaf_243_clk;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire clknet_leaf_242_clk;
 wire _05542_;
 wire _05543_;
 wire clknet_leaf_241_clk;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire clknet_leaf_240_clk;
 wire clknet_leaf_239_clk;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire clknet_leaf_238_clk;
 wire _05571_;
 wire clknet_leaf_237_clk;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire clknet_leaf_236_clk;
 wire _05583_;
 wire clknet_leaf_235_clk;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire clknet_leaf_234_clk;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire clknet_leaf_233_clk;
 wire _05600_;
 wire clknet_leaf_232_clk;
 wire clknet_leaf_231_clk;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire clknet_leaf_230_clk;
 wire _05612_;
 wire _05613_;
 wire clknet_leaf_229_clk;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire clknet_leaf_228_clk;
 wire _05624_;
 wire _05625_;
 wire clknet_leaf_227_clk;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire clknet_leaf_226_clk;
 wire clknet_leaf_225_clk;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire clknet_leaf_224_clk;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire clknet_leaf_223_clk;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire clknet_leaf_222_clk;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_220_clk;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire clknet_leaf_219_clk;
 wire _05690_;
 wire _05691_;
 wire clknet_leaf_218_clk;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire clknet_leaf_217_clk;
 wire _05702_;
 wire _05703_;
 wire clknet_leaf_216_clk;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_214_clk;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire clknet_leaf_213_clk;
 wire _05730_;
 wire clknet_leaf_212_clk;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire clknet_leaf_211_clk;
 wire _05742_;
 wire clknet_leaf_210_clk;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_208_clk;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire clknet_leaf_207_clk;
 wire _05768_;
 wire _05769_;
 wire clknet_leaf_206_clk;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire clknet_leaf_205_clk;
 wire _05780_;
 wire _05781_;
 wire clknet_leaf_204_clk;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_202_clk;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire clknet_leaf_201_clk;
 wire _05808_;
 wire clknet_leaf_200_clk;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire clknet_leaf_199_clk;
 wire _05820_;
 wire clknet_leaf_198_clk;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_196_clk;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire clknet_leaf_195_clk;
 wire _05846_;
 wire _05847_;
 wire clknet_leaf_194_clk;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire clknet_leaf_193_clk;
 wire _05858_;
 wire _05859_;
 wire clknet_leaf_192_clk;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_190_clk;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire clknet_leaf_189_clk;
 wire _05886_;
 wire clknet_leaf_188_clk;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire clknet_leaf_187_clk;
 wire _05898_;
 wire clknet_leaf_186_clk;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_184_clk;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire clknet_leaf_183_clk;
 wire _05924_;
 wire _05925_;
 wire clknet_leaf_182_clk;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire clknet_leaf_181_clk;
 wire _05936_;
 wire _05937_;
 wire clknet_leaf_180_clk;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_178_clk;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire clknet_leaf_177_clk;
 wire _05965_;
 wire clknet_leaf_176_clk;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire clknet_leaf_175_clk;
 wire _05977_;
 wire clknet_leaf_174_clk;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_167_clk;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_163_clk;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire clknet_leaf_160_clk;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire clknet_leaf_159_clk;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire clknet_leaf_156_clk;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire clknet_leaf_152_clk;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire clknet_leaf_150_clk;
 wire _06237_;
 wire clknet_leaf_149_clk;
 wire _06239_;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_146_clk;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_143_clk;
 wire _06275_;
 wire _06276_;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_141_clk;
 wire _06279_;
 wire _06280_;
 wire clknet_leaf_138_clk;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_129_clk;
 wire _06294_;
 wire clknet_leaf_128_clk;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire clknet_leaf_127_clk;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire clknet_leaf_125_clk;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire clknet_leaf_124_clk;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_122_clk;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire clknet_leaf_121_clk;
 wire _06433_;
 wire clknet_leaf_120_clk;
 wire _06435_;
 wire _06436_;
 wire clknet_leaf_119_clk;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire clknet_leaf_117_clk;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire clknet_leaf_116_clk;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire clknet_leaf_115_clk;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire clknet_leaf_114_clk;
 wire _06462_;
 wire _06463_;
 wire clknet_leaf_113_clk;
 wire _06465_;
 wire clknet_leaf_112_clk;
 wire _06467_;
 wire _06468_;
 wire clknet_leaf_110_clk;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire clknet_leaf_109_clk;
 wire _06474_;
 wire _06475_;
 wire clknet_leaf_108_clk;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire clknet_leaf_107_clk;
 wire _06481_;
 wire _06482_;
 wire clknet_leaf_106_clk;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire clknet_leaf_104_clk;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire clknet_leaf_103_clk;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire clknet_leaf_102_clk;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire clknet_leaf_101_clk;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire clknet_leaf_92_clk;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire clknet_leaf_91_clk;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire _06908_;
 wire _06909_;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire clknet_leaf_90_clk;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire clknet_leaf_89_clk;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire clknet_leaf_88_clk;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire clknet_leaf_87_clk;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire clknet_leaf_86_clk;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_82_clk;
 wire _07139_;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_78_clk;
 wire _07144_;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_76_clk;
 wire _07147_;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_73_clk;
 wire _07151_;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_69_clk;
 wire _07156_;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_67_clk;
 wire _07159_;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_65_clk;
 wire _07162_;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_63_clk;
 wire _07165_;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_61_clk;
 wire _07168_;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_59_clk;
 wire _07171_;
 wire clknet_leaf_58_clk;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire clknet_leaf_57_clk;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire clknet_leaf_56_clk;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire clknet_leaf_55_clk;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire clknet_leaf_54_clk;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire clknet_leaf_53_clk;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire clknet_leaf_52_clk;
 wire _07214_;
 wire _07215_;
 wire clknet_leaf_51_clk;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire clknet_leaf_50_clk;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire clknet_leaf_49_clk;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire clknet_leaf_48_clk;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire clknet_leaf_47_clk;
 wire _07242_;
 wire clknet_leaf_46_clk;
 wire _07244_;
 wire clknet_leaf_45_clk;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire clknet_leaf_44_clk;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire clknet_leaf_43_clk;
 wire _07256_;
 wire clknet_leaf_42_clk;
 wire _07258_;
 wire clknet_leaf_41_clk;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire clknet_leaf_40_clk;
 wire _07264_;
 wire clknet_leaf_39_clk;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire clknet_leaf_38_clk;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire clknet_leaf_37_clk;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire clknet_leaf_36_clk;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire clknet_leaf_35_clk;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire clknet_leaf_34_clk;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire clknet_leaf_33_clk;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire clknet_leaf_32_clk;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire clknet_leaf_31_clk;
 wire _07335_;
 wire _07336_;
 wire clknet_leaf_30_clk;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire clknet_leaf_29_clk;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire clknet_leaf_28_clk;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire clknet_leaf_27_clk;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire clknet_leaf_26_clk;
 wire _07363_;
 wire clknet_leaf_25_clk;
 wire _07365_;
 wire clknet_leaf_24_clk;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire clknet_leaf_23_clk;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire clknet_leaf_22_clk;
 wire _07377_;
 wire clknet_leaf_21_clk;
 wire _07379_;
 wire clknet_leaf_20_clk;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire clknet_leaf_19_clk;
 wire _07385_;
 wire clknet_leaf_18_clk;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire clknet_leaf_17_clk;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire _07406_;
 wire _07407_;
 wire _07408_;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire clknet_leaf_16_clk;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire _07420_;
 wire clknet_leaf_15_clk;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire _07436_;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire _07471_;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_11_clk;
 wire _07520_;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_7_clk;
 wire _07525_;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_5_clk;
 wire _07528_;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_2_clk;
 wire _07532_;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_0_clk;
 wire net1039;
 wire net1038;
 wire _07537_;
 wire _07540_;
 wire _07543_;
 wire _07546_;
 wire _07549_;
 wire _07552_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07595_;
 wire _07596_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07623_;
 wire _07625_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07637_;
 wire _07639_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07645_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07716_;
 wire _07717_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07744_;
 wire _07746_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07758_;
 wire _07760_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07766_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire _07932_;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire _07945_;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire _07951_;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire _07980_;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08264_;
 wire _08266_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08283_;
 wire _08284_;
 wire _08288_;
 wire _08289_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08301_;
 wire _08302_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08310_;
 wire _08311_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08374_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire _08444_;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire _08451_;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire _08476_;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08573_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08581_;
 wire _08582_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08599_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08622_;
 wire _08623_;
 wire _08625_;
 wire _08626_;
 wire _08629_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08866_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08905_;
 wire _08940_;
 wire _08944_;
 wire _08948_;
 wire _08952_;
 wire _08956_;
 wire _08960_;
 wire _08965_;
 wire _08969_;
 wire _08973_;
 wire _08977_;
 wire _08981_;
 wire _08985_;
 wire _08989_;
 wire _08993_;
 wire _08997_;
 wire _09001_;
 wire _09005_;
 wire _09009_;
 wire _09014_;
 wire net780;
 wire net779;
 wire net778;
 wire net777;
 wire net776;
 wire net775;
 wire net774;
 wire net773;
 wire net772;
 wire net771;
 wire net770;
 wire net769;
 wire net768;
 wire net767;
 wire net766;
 wire net765;
 wire net764;
 wire net763;
 wire net762;
 wire net761;
 wire net760;
 wire _09050_;
 wire net759;
 wire net758;
 wire net757;
 wire net756;
 wire net755;
 wire net754;
 wire net753;
 wire net752;
 wire net751;
 wire net750;
 wire net749;
 wire net748;
 wire net747;
 wire net746;
 wire net745;
 wire net744;
 wire net743;
 wire net742;
 wire net741;
 wire net740;
 wire net739;
 wire net738;
 wire net737;
 wire net736;
 wire net735;
 wire net734;
 wire net733;
 wire net732;
 wire net731;
 wire net730;
 wire net729;
 wire net728;
 wire net727;
 wire net726;
 wire _09085_;
 wire net725;
 wire net724;
 wire net723;
 wire _09089_;
 wire net722;
 wire net721;
 wire net720;
 wire net719;
 wire _09094_;
 wire net718;
 wire net717;
 wire net716;
 wire _09098_;
 wire net715;
 wire net714;
 wire net713;
 wire _09102_;
 wire net712;
 wire net711;
 wire net710;
 wire _09106_;
 wire net709;
 wire net708;
 wire net707;
 wire _09110_;
 wire net706;
 wire net705;
 wire net704;
 wire _09114_;
 wire net703;
 wire net702;
 wire net701;
 wire _09118_;
 wire net700;
 wire net699;
 wire net698;
 wire _09122_;
 wire net697;
 wire net696;
 wire net695;
 wire _09126_;
 wire net694;
 wire net693;
 wire net692;
 wire _09130_;
 wire net691;
 wire net690;
 wire net689;
 wire _09134_;
 wire net688;
 wire net687;
 wire net686;
 wire _09138_;
 wire net685;
 wire net684;
 wire net683;
 wire _09142_;
 wire net682;
 wire net681;
 wire net680;
 wire _09146_;
 wire net679;
 wire net678;
 wire net677;
 wire _09150_;
 wire net676;
 wire net675;
 wire net674;
 wire _09154_;
 wire net673;
 wire net672;
 wire net671;
 wire net670;
 wire _09159_;
 wire net669;
 wire net668;
 wire net667;
 wire _09163_;
 wire net666;
 wire net665;
 wire net664;
 wire _09167_;
 wire net663;
 wire net662;
 wire net661;
 wire _09171_;
 wire net660;
 wire net659;
 wire net658;
 wire _09175_;
 wire net657;
 wire net656;
 wire net655;
 wire _09179_;
 wire net654;
 wire net653;
 wire net652;
 wire _09183_;
 wire net651;
 wire net650;
 wire net649;
 wire _09187_;
 wire net648;
 wire net647;
 wire net646;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire net645;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire _09290_;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire _09296_;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire _09713_;
 wire net644;
 wire net643;
 wire net642;
 wire net641;
 wire net640;
 wire net639;
 wire net638;
 wire net637;
 wire net636;
 wire net635;
 wire net634;
 wire net633;
 wire _09726_;
 wire _09727_;
 wire net632;
 wire net631;
 wire net630;
 wire _09731_;
 wire net628;
 wire net627;
 wire net626;
 wire _09735_;
 wire _09736_;
 wire net625;
 wire net624;
 wire _09739_;
 wire _09740_;
 wire net623;
 wire _09742_;
 wire net622;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire net621;
 wire net620;
 wire _09755_;
 wire _09756_;
 wire _09757_;
 wire _09758_;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire net619;
 wire _09766_;
 wire _09767_;
 wire net618;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire net617;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire net616;
 wire _09780_;
 wire net615;
 wire net614;
 wire net613;
 wire _09784_;
 wire net612;
 wire _09786_;
 wire _09787_;
 wire net611;
 wire net610;
 wire _09790_;
 wire _09791_;
 wire net609;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire net608;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire net607;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire net606;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire net605;
 wire _09836_;
 wire net604;
 wire _09838_;
 wire net603;
 wire net602;
 wire net601;
 wire net600;
 wire net599;
 wire _09844_;
 wire net598;
 wire net597;
 wire _09847_;
 wire _09848_;
 wire net596;
 wire net595;
 wire net594;
 wire _09852_;
 wire net593;
 wire _09854_;
 wire net592;
 wire _09856_;
 wire _09857_;
 wire net591;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire net590;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire net589;
 wire net588;
 wire _09870_;
 wire net587;
 wire net586;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire net585;
 wire net584;
 wire net583;
 wire _09879_;
 wire net582;
 wire net581;
 wire net580;
 wire net579;
 wire _09884_;
 wire net578;
 wire net577;
 wire _09887_;
 wire net576;
 wire net575;
 wire _09890_;
 wire net574;
 wire net573;
 wire _09893_;
 wire net572;
 wire net571;
 wire _09896_;
 wire net570;
 wire net569;
 wire _09899_;
 wire _09900_;
 wire _09901_;
 wire net568;
 wire net567;
 wire _09904_;
 wire net566;
 wire net565;
 wire net564;
 wire _09908_;
 wire net563;
 wire _09910_;
 wire _09911_;
 wire net562;
 wire _09913_;
 wire net561;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire net560;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire net559;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire net558;
 wire _09936_;
 wire _09937_;
 wire net557;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire net556;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire net555;
 wire _09951_;
 wire _09952_;
 wire _09953_;
 wire net554;
 wire net553;
 wire net552;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire net284;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire net283;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire net282;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire net281;
 wire _09987_;
 wire _09988_;
 wire net280;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire net279;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire net278;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire net277;
 wire net276;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire net275;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire net274;
 wire _10024_;
 wire _10025_;
 wire net273;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire net272;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire net271;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire net270;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire net269;
 wire _10059_;
 wire net268;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire net267;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire net266;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire net265;
 wire _10082_;
 wire _10083_;
 wire net264;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire net263;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire net262;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire net261;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire net260;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire net259;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire net258;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire net257;
 wire _10131_;
 wire _10132_;
 wire net256;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire net255;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire net254;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire net253;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire net252;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire net251;
 wire _10167_;
 wire _10168_;
 wire net250;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire net249;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire net248;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire net247;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire net246;
 wire _10202_;
 wire net245;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire net244;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire net243;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire net242;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire net241;
 wire net240;
 wire net239;
 wire net238;
 wire net237;
 wire net236;
 wire net235;
 wire _10333_;
 wire net234;
 wire net233;
 wire net232;
 wire net231;
 wire _10338_;
 wire net230;
 wire net229;
 wire _10341_;
 wire net228;
 wire net227;
 wire net226;
 wire net225;
 wire _10346_;
 wire net224;
 wire _10348_;
 wire net223;
 wire net222;
 wire _10351_;
 wire _10352_;
 wire net221;
 wire net220;
 wire _10355_;
 wire net219;
 wire net218;
 wire _10358_;
 wire net217;
 wire net216;
 wire _10361_;
 wire net215;
 wire net214;
 wire _10364_;
 wire net213;
 wire net212;
 wire _10367_;
 wire net211;
 wire net210;
 wire net209;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire net208;
 wire net207;
 wire net206;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire net205;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire net204;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire net203;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire net202;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire net201;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire net200;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire net199;
 wire _10434_;
 wire _10435_;
 wire _10436_;
 wire _10437_;
 wire net198;
 wire _10439_;
 wire _10440_;
 wire net197;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire net196;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire net195;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire _10454_;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire net194;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire net193;
 wire _10463_;
 wire _10464_;
 wire net192;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire net191;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire net190;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire net189;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire net188;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire net187;
 wire net186;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire net185;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire net184;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire net183;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire net182;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire net181;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire net180;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire net179;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire net178;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire net177;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire net176;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire net175;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire net174;
 wire _10583_;
 wire _10584_;
 wire net173;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire net172;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire net171;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire net170;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire net169;
 wire _10607_;
 wire _10608_;
 wire net168;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire net167;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire net166;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire net165;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire net164;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire net163;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire net162;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire net161;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire net160;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire net159;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire net158;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire _10676_;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire net157;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire net156;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire net155;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire net154;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire net153;
 wire net152;
 wire net151;
 wire net150;
 wire net149;
 wire net148;
 wire net147;
 wire net146;
 wire net145;
 wire _10812_;
 wire net144;
 wire net143;
 wire net142;
 wire net141;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire net140;
 wire net139;
 wire net138;
 wire net137;
 wire net136;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire net135;
 wire net134;
 wire _10833_;
 wire net133;
 wire net132;
 wire net131;
 wire _10837_;
 wire net130;
 wire net129;
 wire _10840_;
 wire net128;
 wire net127;
 wire _10843_;
 wire net126;
 wire net125;
 wire _10846_;
 wire net124;
 wire net123;
 wire _10849_;
 wire net122;
 wire _10851_;
 wire net121;
 wire net120;
 wire _10854_;
 wire net119;
 wire net118;
 wire _10857_;
 wire net117;
 wire net116;
 wire _10860_;
 wire net115;
 wire net114;
 wire _10863_;
 wire net113;
 wire _10865_;
 wire net112;
 wire net111;
 wire _10868_;
 wire net110;
 wire net109;
 wire _10871_;
 wire net108;
 wire _10873_;
 wire net107;
 wire _10875_;
 wire net106;
 wire net105;
 wire _10878_;
 wire net104;
 wire net103;
 wire _10881_;
 wire net102;
 wire net101;
 wire _10884_;
 wire net100;
 wire _10886_;
 wire net99;
 wire net98;
 wire _10889_;
 wire net97;
 wire net96;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire net95;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire net94;
 wire net93;
 wire net92;
 wire net91;
 wire net90;
 wire net89;
 wire net88;
 wire net87;
 wire net86;
 wire net85;
 wire _10940_;
 wire net84;
 wire net83;
 wire _10943_;
 wire _10944_;
 wire net82;
 wire net81;
 wire _10947_;
 wire net80;
 wire net79;
 wire net78;
 wire net77;
 wire net76;
 wire _10953_;
 wire _10954_;
 wire net75;
 wire net74;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire net73;
 wire net72;
 wire _10963_;
 wire net71;
 wire net70;
 wire net69;
 wire _10967_;
 wire net68;
 wire net67;
 wire _10970_;
 wire net66;
 wire net65;
 wire _10973_;
 wire net64;
 wire net63;
 wire _10976_;
 wire net62;
 wire net61;
 wire _10979_;
 wire net60;
 wire net59;
 wire _10982_;
 wire net58;
 wire _10984_;
 wire net57;
 wire net56;
 wire _10987_;
 wire net55;
 wire net54;
 wire _10990_;
 wire net53;
 wire net52;
 wire _10993_;
 wire net51;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire net50;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire net49;
 wire _11017_;
 wire net48;
 wire net47;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire net46;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire net45;
 wire _11059_;
 wire _11060_;
 wire net44;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire net43;
 wire _11070_;
 wire _11071_;
 wire net42;
 wire _11073_;
 wire net41;
 wire _11075_;
 wire _11076_;
 wire net40;
 wire net39;
 wire _11079_;
 wire net38;
 wire net37;
 wire _11082_;
 wire _11083_;
 wire net36;
 wire net35;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire net34;
 wire net33;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire net32;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire net31;
 wire _11116_;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire net30;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire net29;
 wire _11132_;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire net28;
 wire net27;
 wire _11140_;
 wire _11141_;
 wire net26;
 wire _11143_;
 wire net25;
 wire _11145_;
 wire net24;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire _11165_;
 wire net23;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire net22;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire net21;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire _11213_;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire net20;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire _11302_;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire _11311_;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire net19;
 wire net18;
 wire _11515_;
 wire net17;
 wire net16;
 wire _11518_;
 wire net15;
 wire net14;
 wire _11521_;
 wire net13;
 wire net12;
 wire _11524_;
 wire net11;
 wire net10;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire net9;
 wire net8;
 wire _11532_;
 wire net7;
 wire net6;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire net5;
 wire net4;
 wire _11541_;
 wire net3;
 wire net2;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire _11854_;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire _11935_;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire _12048_;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire _12507_;
 wire _12508_;
 wire _12509_;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire _12528_;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire _12585_;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire clknet_leaf_126_clk;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire _12641_;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire _12648_;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire _12653_;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire _12671_;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire clknet_leaf_93_clk;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire _13239_;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire _13312_;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire _13318_;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire _13388_;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire clknet_leaf_134_clk;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire _13841_;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire _13955_;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire _13979_;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire \count15_1[1] ;
 wire \count15_1[2] ;
 wire \count15_1[3] ;
 wire \count15_1[4] ;
 wire \count15_1[5] ;
 wire \count15_2[1] ;
 wire \count15_2[2] ;
 wire \count15_2[3] ;
 wire \count15_2[4] ;
 wire \count15_2[5] ;
 wire \count16_1[1] ;
 wire \count16_1[2] ;
 wire \count16_1[3] ;
 wire \count16_1[4] ;
 wire \count16_1[5] ;
 wire \count16_2[1] ;
 wire \count16_2[2] ;
 wire \count16_2[3] ;
 wire \count16_2[4] ;
 wire \count16_2[5] ;
 wire \count2_1[1] ;
 wire \count2_1[2] ;
 wire \count2_1[3] ;
 wire \count2_1[4] ;
 wire \count2_1[5] ;
 wire \count2_2[1] ;
 wire \count2_2[2] ;
 wire \count2_2[3] ;
 wire \count2_2[4] ;
 wire \count2_2[5] ;
 wire \count7_1[1] ;
 wire \count7_1[2] ;
 wire \count7_1[3] ;
 wire \count7_1[4] ;
 wire \count7_1[5] ;
 wire \count7_2[1] ;
 wire \count7_2[2] ;
 wire \count7_2[3] ;
 wire \count7_2[4] ;
 wire \count7_2[5] ;
 wire \count_1[1] ;
 wire \count_1[2] ;
 wire \count_1[3] ;
 wire \count_1[4] ;
 wire \count_1[5] ;
 wire \count_2[1] ;
 wire \count_2[2] ;
 wire \count_2[3] ;
 wire \count_2[4] ;
 wire \count_2[5] ;
 wire \count_2[6] ;
 wire \count_hash1[1] ;
 wire \count_hash1[2] ;
 wire \count_hash1[3] ;
 wire \count_hash1[4] ;
 wire \count_hash1[5] ;
 wire \count_hash1[6] ;
 wire \count_hash2[1] ;
 wire \count_hash2[2] ;
 wire \count_hash2[3] ;
 wire \count_hash2[4] ;
 wire \count_hash2[5] ;
 wire done;
 wire \hash.CA1.S0.X[0] ;
 wire \hash.CA1.S0.X[10] ;
 wire \hash.CA1.S0.X[11] ;
 wire \hash.CA1.S0.X[12] ;
 wire \hash.CA1.S0.X[13] ;
 wire \hash.CA1.S0.X[14] ;
 wire \hash.CA1.S0.X[15] ;
 wire \hash.CA1.S0.X[16] ;
 wire \hash.CA1.S0.X[17] ;
 wire \hash.CA1.S0.X[18] ;
 wire \hash.CA1.S0.X[19] ;
 wire \hash.CA1.S0.X[1] ;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_157_clk;
 wire \hash.CA1.S0.X[22] ;
 wire \hash.CA1.S0.X[23] ;
 wire clknet_leaf_155_clk;
 wire \hash.CA1.S0.X[25] ;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_153_clk;
 wire \hash.CA1.S0.X[28] ;
 wire \hash.CA1.S0.X[29] ;
 wire \hash.CA1.S0.X[2] ;
 wire clknet_leaf_151_clk;
 wire \hash.CA1.S0.X[31] ;
 wire \hash.CA1.S0.X[3] ;
 wire clknet_leaf_162_clk;
 wire \hash.CA1.S0.X[5] ;
 wire \hash.CA1.S0.X[6] ;
 wire \hash.CA1.S0.X[7] ;
 wire clknet_leaf_161_clk;
 wire \hash.CA1.S0.X[9] ;
 wire \hash.CA1.S1.X[0] ;
 wire \hash.CA1.S1.X[10] ;
 wire clknet_leaf_99_clk;
 wire \hash.CA1.S1.X[12] ;
 wire \hash.CA1.S1.X[13] ;
 wire \hash.CA1.S1.X[14] ;
 wire clknet_leaf_98_clk;
 wire \hash.CA1.S1.X[16] ;
 wire \hash.CA1.S1.X[17] ;
 wire \hash.CA1.S1.X[18] ;
 wire \hash.CA1.S1.X[19] ;
 wire \hash.CA1.S1.X[1] ;
 wire \hash.CA1.S1.X[20] ;
 wire \hash.CA1.S1.X[21] ;
 wire \hash.CA1.S1.X[22] ;
 wire \hash.CA1.S1.X[23] ;
 wire \hash.CA1.S1.X[24] ;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_94_clk;
 wire \hash.CA1.S1.X[29] ;
 wire \hash.CA1.S1.X[2] ;
 wire \hash.CA1.S1.X[30] ;
 wire \hash.CA1.S1.X[31] ;
 wire \hash.CA1.S1.X[3] ;
 wire \hash.CA1.S1.X[4] ;
 wire \hash.CA1.S1.X[5] ;
 wire \hash.CA1.S1.X[6] ;
 wire \hash.CA1.S1.X[7] ;
 wire clknet_leaf_100_clk;
 wire \hash.CA1.S1.X[9] ;
 wire \hash.CA1.b[0] ;
 wire \hash.CA1.b[10] ;
 wire \hash.CA1.b[11] ;
 wire clknet_leaf_137_clk;
 wire \hash.CA1.b[13] ;
 wire \hash.CA1.b[14] ;
 wire \hash.CA1.b[15] ;
 wire \hash.CA1.b[16] ;
 wire \hash.CA1.b[17] ;
 wire \hash.CA1.b[18] ;
 wire clknet_leaf_136_clk;
 wire \hash.CA1.b[1] ;
 wire \hash.CA1.b[20] ;
 wire \hash.CA1.b[21] ;
 wire \hash.CA1.b[22] ;
 wire clknet_leaf_135_clk;
 wire \hash.CA1.b[24] ;
 wire \hash.CA1.b[25] ;
 wire \hash.CA1.b[26] ;
 wire \hash.CA1.b[27] ;
 wire \hash.CA1.b[28] ;
 wire \hash.CA1.b[29] ;
 wire \hash.CA1.b[2] ;
 wire \hash.CA1.b[30] ;
 wire \hash.CA1.b[31] ;
 wire \hash.CA1.b[3] ;
 wire \hash.CA1.b[4] ;
 wire \hash.CA1.b[5] ;
 wire \hash.CA1.b[6] ;
 wire \hash.CA1.b[7] ;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_139_clk;
 wire \hash.CA1.c[0] ;
 wire \hash.CA1.d[0] ;
 wire \hash.CA1.f[0] ;
 wire \hash.CA1.f[10] ;
 wire \hash.CA1.f[11] ;
 wire \hash.CA1.f[12] ;
 wire \hash.CA1.f[13] ;
 wire \hash.CA1.f[14] ;
 wire \hash.CA1.f[15] ;
 wire \hash.CA1.f[16] ;
 wire \hash.CA1.f[17] ;
 wire clknet_leaf_111_clk;
 wire \hash.CA1.f[19] ;
 wire \hash.CA1.f[1] ;
 wire \hash.CA1.f[20] ;
 wire \hash.CA1.f[21] ;
 wire \hash.CA1.f[22] ;
 wire \hash.CA1.f[23] ;
 wire clknet_leaf_105_clk;
 wire \hash.CA1.f[25] ;
 wire \hash.CA1.f[26] ;
 wire \hash.CA1.f[27] ;
 wire \hash.CA1.f[28] ;
 wire \hash.CA1.f[29] ;
 wire \hash.CA1.f[2] ;
 wire \hash.CA1.f[30] ;
 wire \hash.CA1.f[31] ;
 wire \hash.CA1.f[3] ;
 wire \hash.CA1.f[4] ;
 wire \hash.CA1.f[5] ;
 wire \hash.CA1.f[6] ;
 wire \hash.CA1.f[7] ;
 wire \hash.CA1.f[8] ;
 wire clknet_leaf_118_clk;
 wire \hash.CA1.k_i1[0] ;
 wire \hash.CA1.k_i1[10] ;
 wire \hash.CA1.k_i1[11] ;
 wire \hash.CA1.k_i1[12] ;
 wire \hash.CA1.k_i1[13] ;
 wire \hash.CA1.k_i1[14] ;
 wire \hash.CA1.k_i1[15] ;
 wire \hash.CA1.k_i1[16] ;
 wire \hash.CA1.k_i1[17] ;
 wire \hash.CA1.k_i1[18] ;
 wire \hash.CA1.k_i1[19] ;
 wire \hash.CA1.k_i1[1] ;
 wire \hash.CA1.k_i1[20] ;
 wire \hash.CA1.k_i1[21] ;
 wire \hash.CA1.k_i1[22] ;
 wire \hash.CA1.k_i1[23] ;
 wire \hash.CA1.k_i1[24] ;
 wire \hash.CA1.k_i1[25] ;
 wire \hash.CA1.k_i1[26] ;
 wire \hash.CA1.k_i1[27] ;
 wire \hash.CA1.k_i1[28] ;
 wire \hash.CA1.k_i1[29] ;
 wire \hash.CA1.k_i1[2] ;
 wire \hash.CA1.k_i1[30] ;
 wire \hash.CA1.k_i1[31] ;
 wire \hash.CA1.k_i1[3] ;
 wire \hash.CA1.k_i1[4] ;
 wire \hash.CA1.k_i1[5] ;
 wire \hash.CA1.k_i1[6] ;
 wire \hash.CA1.k_i1[7] ;
 wire \hash.CA1.k_i1[8] ;
 wire \hash.CA1.k_i1[9] ;
 wire \hash.CA1.k_i2[0] ;
 wire \hash.CA1.k_i2[10] ;
 wire \hash.CA1.k_i2[11] ;
 wire \hash.CA1.k_i2[12] ;
 wire \hash.CA1.k_i2[13] ;
 wire \hash.CA1.k_i2[14] ;
 wire \hash.CA1.k_i2[15] ;
 wire \hash.CA1.k_i2[16] ;
 wire \hash.CA1.k_i2[17] ;
 wire \hash.CA1.k_i2[18] ;
 wire \hash.CA1.k_i2[19] ;
 wire \hash.CA1.k_i2[1] ;
 wire \hash.CA1.k_i2[20] ;
 wire \hash.CA1.k_i2[21] ;
 wire \hash.CA1.k_i2[22] ;
 wire \hash.CA1.k_i2[23] ;
 wire \hash.CA1.k_i2[24] ;
 wire \hash.CA1.k_i2[25] ;
 wire \hash.CA1.k_i2[26] ;
 wire \hash.CA1.k_i2[27] ;
 wire \hash.CA1.k_i2[28] ;
 wire \hash.CA1.k_i2[29] ;
 wire \hash.CA1.k_i2[2] ;
 wire \hash.CA1.k_i2[30] ;
 wire \hash.CA1.k_i2[31] ;
 wire \hash.CA1.k_i2[3] ;
 wire \hash.CA1.k_i2[4] ;
 wire \hash.CA1.k_i2[5] ;
 wire \hash.CA1.k_i2[6] ;
 wire \hash.CA1.k_i2[7] ;
 wire \hash.CA1.k_i2[8] ;
 wire \hash.CA1.k_i2[9] ;
 wire \hash.CA1.p1[0] ;
 wire \hash.CA1.p1[10] ;
 wire \hash.CA1.p1[11] ;
 wire \hash.CA1.p1[12] ;
 wire \hash.CA1.p1[13] ;
 wire \hash.CA1.p1[14] ;
 wire \hash.CA1.p1[15] ;
 wire \hash.CA1.p1[16] ;
 wire \hash.CA1.p1[17] ;
 wire \hash.CA1.p1[18] ;
 wire \hash.CA1.p1[19] ;
 wire \hash.CA1.p1[1] ;
 wire \hash.CA1.p1[20] ;
 wire \hash.CA1.p1[21] ;
 wire \hash.CA1.p1[22] ;
 wire \hash.CA1.p1[23] ;
 wire \hash.CA1.p1[24] ;
 wire \hash.CA1.p1[25] ;
 wire \hash.CA1.p1[26] ;
 wire \hash.CA1.p1[27] ;
 wire \hash.CA1.p1[28] ;
 wire \hash.CA1.p1[29] ;
 wire \hash.CA1.p1[2] ;
 wire \hash.CA1.p1[30] ;
 wire \hash.CA1.p1[31] ;
 wire \hash.CA1.p1[3] ;
 wire \hash.CA1.p1[4] ;
 wire \hash.CA1.p1[5] ;
 wire \hash.CA1.p1[6] ;
 wire \hash.CA1.p1[7] ;
 wire \hash.CA1.p1[8] ;
 wire \hash.CA1.p1[9] ;
 wire \hash.CA1.p2[0] ;
 wire \hash.CA1.p2[10] ;
 wire \hash.CA1.p2[11] ;
 wire \hash.CA1.p2[12] ;
 wire \hash.CA1.p2[13] ;
 wire \hash.CA1.p2[14] ;
 wire \hash.CA1.p2[15] ;
 wire \hash.CA1.p2[16] ;
 wire \hash.CA1.p2[17] ;
 wire \hash.CA1.p2[18] ;
 wire \hash.CA1.p2[19] ;
 wire \hash.CA1.p2[1] ;
 wire \hash.CA1.p2[20] ;
 wire \hash.CA1.p2[21] ;
 wire \hash.CA1.p2[22] ;
 wire \hash.CA1.p2[23] ;
 wire \hash.CA1.p2[24] ;
 wire \hash.CA1.p2[25] ;
 wire \hash.CA1.p2[26] ;
 wire \hash.CA1.p2[27] ;
 wire \hash.CA1.p2[28] ;
 wire \hash.CA1.p2[29] ;
 wire \hash.CA1.p2[2] ;
 wire \hash.CA1.p2[30] ;
 wire \hash.CA1.p2[31] ;
 wire \hash.CA1.p2[3] ;
 wire \hash.CA1.p2[4] ;
 wire \hash.CA1.p2[5] ;
 wire \hash.CA1.p2[6] ;
 wire \hash.CA1.p2[7] ;
 wire \hash.CA1.p2[8] ;
 wire \hash.CA1.p2[9] ;
 wire \hash.CA1.p3[0] ;
 wire \hash.CA1.p3[10] ;
 wire \hash.CA1.p3[11] ;
 wire \hash.CA1.p3[12] ;
 wire \hash.CA1.p3[13] ;
 wire \hash.CA1.p3[14] ;
 wire \hash.CA1.p3[15] ;
 wire \hash.CA1.p3[16] ;
 wire \hash.CA1.p3[17] ;
 wire \hash.CA1.p3[18] ;
 wire \hash.CA1.p3[19] ;
 wire \hash.CA1.p3[1] ;
 wire \hash.CA1.p3[20] ;
 wire \hash.CA1.p3[21] ;
 wire \hash.CA1.p3[22] ;
 wire \hash.CA1.p3[23] ;
 wire \hash.CA1.p3[24] ;
 wire \hash.CA1.p3[25] ;
 wire \hash.CA1.p3[26] ;
 wire \hash.CA1.p3[27] ;
 wire \hash.CA1.p3[28] ;
 wire \hash.CA1.p3[29] ;
 wire \hash.CA1.p3[2] ;
 wire \hash.CA1.p3[30] ;
 wire \hash.CA1.p3[31] ;
 wire \hash.CA1.p3[3] ;
 wire \hash.CA1.p3[4] ;
 wire \hash.CA1.p3[5] ;
 wire \hash.CA1.p3[6] ;
 wire \hash.CA1.p3[7] ;
 wire \hash.CA1.p3[8] ;
 wire \hash.CA1.p3[9] ;
 wire \hash.CA1.p4[0] ;
 wire \hash.CA1.p4[10] ;
 wire \hash.CA1.p4[11] ;
 wire \hash.CA1.p4[12] ;
 wire \hash.CA1.p4[13] ;
 wire \hash.CA1.p4[14] ;
 wire \hash.CA1.p4[15] ;
 wire \hash.CA1.p4[16] ;
 wire \hash.CA1.p4[17] ;
 wire \hash.CA1.p4[18] ;
 wire \hash.CA1.p4[19] ;
 wire \hash.CA1.p4[1] ;
 wire \hash.CA1.p4[20] ;
 wire \hash.CA1.p4[21] ;
 wire \hash.CA1.p4[22] ;
 wire \hash.CA1.p4[23] ;
 wire \hash.CA1.p4[24] ;
 wire \hash.CA1.p4[25] ;
 wire \hash.CA1.p4[26] ;
 wire \hash.CA1.p4[27] ;
 wire \hash.CA1.p4[28] ;
 wire \hash.CA1.p4[29] ;
 wire \hash.CA1.p4[2] ;
 wire \hash.CA1.p4[30] ;
 wire \hash.CA1.p4[31] ;
 wire \hash.CA1.p4[3] ;
 wire \hash.CA1.p4[4] ;
 wire \hash.CA1.p4[5] ;
 wire \hash.CA1.p4[6] ;
 wire \hash.CA1.p4[7] ;
 wire \hash.CA1.p4[8] ;
 wire \hash.CA1.p4[9] ;
 wire \hash.CA1.p5[0] ;
 wire \hash.CA1.p5[10] ;
 wire \hash.CA1.p5[11] ;
 wire \hash.CA1.p5[12] ;
 wire \hash.CA1.p5[13] ;
 wire \hash.CA1.p5[14] ;
 wire \hash.CA1.p5[15] ;
 wire \hash.CA1.p5[16] ;
 wire \hash.CA1.p5[17] ;
 wire \hash.CA1.p5[18] ;
 wire \hash.CA1.p5[19] ;
 wire \hash.CA1.p5[1] ;
 wire \hash.CA1.p5[20] ;
 wire \hash.CA1.p5[21] ;
 wire \hash.CA1.p5[22] ;
 wire \hash.CA1.p5[23] ;
 wire \hash.CA1.p5[24] ;
 wire \hash.CA1.p5[25] ;
 wire \hash.CA1.p5[26] ;
 wire \hash.CA1.p5[27] ;
 wire \hash.CA1.p5[28] ;
 wire \hash.CA1.p5[29] ;
 wire \hash.CA1.p5[2] ;
 wire \hash.CA1.p5[30] ;
 wire \hash.CA1.p5[31] ;
 wire \hash.CA1.p5[3] ;
 wire \hash.CA1.p5[4] ;
 wire \hash.CA1.p5[5] ;
 wire \hash.CA1.p5[6] ;
 wire \hash.CA1.p5[7] ;
 wire \hash.CA1.p5[8] ;
 wire \hash.CA1.p5[9] ;
 wire \hash.CA1.w_i1[0] ;
 wire \hash.CA1.w_i1[10] ;
 wire \hash.CA1.w_i1[11] ;
 wire \hash.CA1.w_i1[12] ;
 wire \hash.CA1.w_i1[13] ;
 wire \hash.CA1.w_i1[14] ;
 wire \hash.CA1.w_i1[15] ;
 wire \hash.CA1.w_i1[16] ;
 wire \hash.CA1.w_i1[17] ;
 wire \hash.CA1.w_i1[18] ;
 wire \hash.CA1.w_i1[19] ;
 wire \hash.CA1.w_i1[1] ;
 wire \hash.CA1.w_i1[20] ;
 wire \hash.CA1.w_i1[21] ;
 wire \hash.CA1.w_i1[22] ;
 wire \hash.CA1.w_i1[23] ;
 wire \hash.CA1.w_i1[24] ;
 wire \hash.CA1.w_i1[25] ;
 wire \hash.CA1.w_i1[26] ;
 wire \hash.CA1.w_i1[27] ;
 wire \hash.CA1.w_i1[28] ;
 wire \hash.CA1.w_i1[29] ;
 wire \hash.CA1.w_i1[2] ;
 wire \hash.CA1.w_i1[30] ;
 wire \hash.CA1.w_i1[31] ;
 wire \hash.CA1.w_i1[3] ;
 wire \hash.CA1.w_i1[4] ;
 wire \hash.CA1.w_i1[5] ;
 wire \hash.CA1.w_i1[6] ;
 wire \hash.CA1.w_i1[7] ;
 wire \hash.CA1.w_i1[8] ;
 wire \hash.CA1.w_i1[9] ;
 wire \hash.CA1.w_i2[0] ;
 wire \hash.CA1.w_i2[10] ;
 wire \hash.CA1.w_i2[11] ;
 wire \hash.CA1.w_i2[12] ;
 wire \hash.CA1.w_i2[13] ;
 wire \hash.CA1.w_i2[14] ;
 wire \hash.CA1.w_i2[15] ;
 wire \hash.CA1.w_i2[16] ;
 wire \hash.CA1.w_i2[17] ;
 wire \hash.CA1.w_i2[18] ;
 wire \hash.CA1.w_i2[19] ;
 wire \hash.CA1.w_i2[1] ;
 wire \hash.CA1.w_i2[20] ;
 wire \hash.CA1.w_i2[21] ;
 wire \hash.CA1.w_i2[22] ;
 wire \hash.CA1.w_i2[23] ;
 wire \hash.CA1.w_i2[24] ;
 wire \hash.CA1.w_i2[25] ;
 wire \hash.CA1.w_i2[26] ;
 wire \hash.CA1.w_i2[27] ;
 wire \hash.CA1.w_i2[28] ;
 wire \hash.CA1.w_i2[29] ;
 wire \hash.CA1.w_i2[2] ;
 wire \hash.CA1.w_i2[30] ;
 wire \hash.CA1.w_i2[31] ;
 wire \hash.CA1.w_i2[3] ;
 wire \hash.CA1.w_i2[4] ;
 wire \hash.CA1.w_i2[5] ;
 wire \hash.CA1.w_i2[6] ;
 wire \hash.CA1.w_i2[7] ;
 wire \hash.CA1.w_i2[8] ;
 wire \hash.CA1.w_i2[9] ;
 wire \hash.CA2.S1.X[0] ;
 wire \hash.CA2.S1.X[10] ;
 wire \hash.CA2.S1.X[11] ;
 wire \hash.CA2.S1.X[12] ;
 wire \hash.CA2.S1.X[13] ;
 wire \hash.CA2.S1.X[14] ;
 wire \hash.CA2.S1.X[15] ;
 wire \hash.CA2.S1.X[16] ;
 wire \hash.CA2.S1.X[17] ;
 wire \hash.CA2.S1.X[18] ;
 wire \hash.CA2.S1.X[19] ;
 wire \hash.CA2.S1.X[1] ;
 wire \hash.CA2.S1.X[20] ;
 wire \hash.CA2.S1.X[21] ;
 wire \hash.CA2.S1.X[22] ;
 wire \hash.CA2.S1.X[23] ;
 wire \hash.CA2.S1.X[24] ;
 wire \hash.CA2.S1.X[25] ;
 wire \hash.CA2.S1.X[26] ;
 wire \hash.CA2.S1.X[27] ;
 wire \hash.CA2.S1.X[28] ;
 wire \hash.CA2.S1.X[29] ;
 wire \hash.CA2.S1.X[2] ;
 wire \hash.CA2.S1.X[30] ;
 wire \hash.CA2.S1.X[31] ;
 wire \hash.CA2.S1.X[3] ;
 wire \hash.CA2.S1.X[4] ;
 wire \hash.CA2.S1.X[5] ;
 wire \hash.CA2.S1.X[6] ;
 wire \hash.CA2.S1.X[7] ;
 wire \hash.CA2.S1.X[8] ;
 wire \hash.CA2.S1.X[9] ;
 wire \hash.CA2.a_dash[0] ;
 wire \hash.CA2.a_dash[10] ;
 wire \hash.CA2.a_dash[11] ;
 wire \hash.CA2.a_dash[12] ;
 wire \hash.CA2.a_dash[13] ;
 wire \hash.CA2.a_dash[14] ;
 wire \hash.CA2.a_dash[15] ;
 wire \hash.CA2.a_dash[16] ;
 wire \hash.CA2.a_dash[17] ;
 wire \hash.CA2.a_dash[18] ;
 wire \hash.CA2.a_dash[19] ;
 wire \hash.CA2.a_dash[1] ;
 wire \hash.CA2.a_dash[20] ;
 wire \hash.CA2.a_dash[21] ;
 wire \hash.CA2.a_dash[22] ;
 wire \hash.CA2.a_dash[23] ;
 wire \hash.CA2.a_dash[24] ;
 wire \hash.CA2.a_dash[25] ;
 wire \hash.CA2.a_dash[26] ;
 wire \hash.CA2.a_dash[27] ;
 wire \hash.CA2.a_dash[28] ;
 wire \hash.CA2.a_dash[29] ;
 wire \hash.CA2.a_dash[2] ;
 wire \hash.CA2.a_dash[30] ;
 wire \hash.CA2.a_dash[31] ;
 wire \hash.CA2.a_dash[3] ;
 wire \hash.CA2.a_dash[4] ;
 wire \hash.CA2.a_dash[5] ;
 wire \hash.CA2.a_dash[6] ;
 wire \hash.CA2.a_dash[7] ;
 wire \hash.CA2.a_dash[8] ;
 wire \hash.CA2.a_dash[9] ;
 wire \hash.CA2.b_dash[0] ;
 wire \hash.CA2.b_dash[10] ;
 wire \hash.CA2.b_dash[11] ;
 wire \hash.CA2.b_dash[12] ;
 wire \hash.CA2.b_dash[13] ;
 wire \hash.CA2.b_dash[14] ;
 wire \hash.CA2.b_dash[15] ;
 wire \hash.CA2.b_dash[16] ;
 wire \hash.CA2.b_dash[17] ;
 wire \hash.CA2.b_dash[18] ;
 wire \hash.CA2.b_dash[19] ;
 wire \hash.CA2.b_dash[1] ;
 wire \hash.CA2.b_dash[20] ;
 wire \hash.CA2.b_dash[21] ;
 wire \hash.CA2.b_dash[22] ;
 wire \hash.CA2.b_dash[23] ;
 wire \hash.CA2.b_dash[24] ;
 wire \hash.CA2.b_dash[25] ;
 wire \hash.CA2.b_dash[26] ;
 wire \hash.CA2.b_dash[27] ;
 wire \hash.CA2.b_dash[28] ;
 wire \hash.CA2.b_dash[29] ;
 wire \hash.CA2.b_dash[2] ;
 wire \hash.CA2.b_dash[30] ;
 wire \hash.CA2.b_dash[31] ;
 wire \hash.CA2.b_dash[3] ;
 wire \hash.CA2.b_dash[4] ;
 wire \hash.CA2.b_dash[5] ;
 wire \hash.CA2.b_dash[6] ;
 wire \hash.CA2.b_dash[7] ;
 wire \hash.CA2.b_dash[8] ;
 wire \hash.CA2.b_dash[9] ;
 wire \hash.CA2.e_dash[0] ;
 wire \hash.CA2.e_dash[10] ;
 wire \hash.CA2.e_dash[11] ;
 wire \hash.CA2.e_dash[12] ;
 wire \hash.CA2.e_dash[13] ;
 wire \hash.CA2.e_dash[14] ;
 wire \hash.CA2.e_dash[15] ;
 wire \hash.CA2.e_dash[16] ;
 wire \hash.CA2.e_dash[17] ;
 wire \hash.CA2.e_dash[18] ;
 wire \hash.CA2.e_dash[19] ;
 wire \hash.CA2.e_dash[1] ;
 wire \hash.CA2.e_dash[20] ;
 wire \hash.CA2.e_dash[21] ;
 wire \hash.CA2.e_dash[22] ;
 wire \hash.CA2.e_dash[23] ;
 wire \hash.CA2.e_dash[24] ;
 wire \hash.CA2.e_dash[25] ;
 wire \hash.CA2.e_dash[26] ;
 wire \hash.CA2.e_dash[27] ;
 wire \hash.CA2.e_dash[28] ;
 wire \hash.CA2.e_dash[29] ;
 wire \hash.CA2.e_dash[2] ;
 wire \hash.CA2.e_dash[30] ;
 wire \hash.CA2.e_dash[31] ;
 wire \hash.CA2.e_dash[3] ;
 wire \hash.CA2.e_dash[4] ;
 wire \hash.CA2.e_dash[5] ;
 wire \hash.CA2.e_dash[6] ;
 wire \hash.CA2.e_dash[7] ;
 wire \hash.CA2.e_dash[8] ;
 wire \hash.CA2.e_dash[9] ;
 wire \hash.CA2.f_dash[0] ;
 wire \hash.CA2.f_dash[10] ;
 wire \hash.CA2.f_dash[11] ;
 wire \hash.CA2.f_dash[12] ;
 wire \hash.CA2.f_dash[13] ;
 wire \hash.CA2.f_dash[14] ;
 wire \hash.CA2.f_dash[15] ;
 wire \hash.CA2.f_dash[16] ;
 wire \hash.CA2.f_dash[17] ;
 wire \hash.CA2.f_dash[18] ;
 wire \hash.CA2.f_dash[19] ;
 wire \hash.CA2.f_dash[1] ;
 wire \hash.CA2.f_dash[20] ;
 wire \hash.CA2.f_dash[21] ;
 wire \hash.CA2.f_dash[22] ;
 wire \hash.CA2.f_dash[23] ;
 wire \hash.CA2.f_dash[24] ;
 wire \hash.CA2.f_dash[25] ;
 wire \hash.CA2.f_dash[26] ;
 wire \hash.CA2.f_dash[27] ;
 wire \hash.CA2.f_dash[28] ;
 wire \hash.CA2.f_dash[29] ;
 wire \hash.CA2.f_dash[2] ;
 wire \hash.CA2.f_dash[30] ;
 wire \hash.CA2.f_dash[31] ;
 wire \hash.CA2.f_dash[3] ;
 wire \hash.CA2.f_dash[4] ;
 wire \hash.CA2.f_dash[5] ;
 wire \hash.CA2.f_dash[6] ;
 wire \hash.CA2.f_dash[7] ;
 wire \hash.CA2.f_dash[8] ;
 wire \hash.CA2.f_dash[9] ;
 wire \hash.CA2.p1[0] ;
 wire \hash.CA2.p1[10] ;
 wire \hash.CA2.p1[11] ;
 wire \hash.CA2.p1[12] ;
 wire \hash.CA2.p1[13] ;
 wire \hash.CA2.p1[14] ;
 wire \hash.CA2.p1[15] ;
 wire \hash.CA2.p1[16] ;
 wire \hash.CA2.p1[17] ;
 wire \hash.CA2.p1[18] ;
 wire \hash.CA2.p1[19] ;
 wire \hash.CA2.p1[1] ;
 wire \hash.CA2.p1[20] ;
 wire \hash.CA2.p1[21] ;
 wire \hash.CA2.p1[22] ;
 wire \hash.CA2.p1[23] ;
 wire \hash.CA2.p1[24] ;
 wire \hash.CA2.p1[25] ;
 wire \hash.CA2.p1[26] ;
 wire \hash.CA2.p1[27] ;
 wire \hash.CA2.p1[28] ;
 wire \hash.CA2.p1[29] ;
 wire \hash.CA2.p1[2] ;
 wire \hash.CA2.p1[30] ;
 wire \hash.CA2.p1[31] ;
 wire \hash.CA2.p1[3] ;
 wire \hash.CA2.p1[4] ;
 wire \hash.CA2.p1[5] ;
 wire \hash.CA2.p1[6] ;
 wire \hash.CA2.p1[7] ;
 wire \hash.CA2.p1[8] ;
 wire \hash.CA2.p1[9] ;
 wire \hash.CA2.p3[0] ;
 wire \hash.CA2.p3[10] ;
 wire \hash.CA2.p3[11] ;
 wire \hash.CA2.p3[12] ;
 wire \hash.CA2.p3[13] ;
 wire \hash.CA2.p3[14] ;
 wire \hash.CA2.p3[15] ;
 wire \hash.CA2.p3[16] ;
 wire \hash.CA2.p3[17] ;
 wire \hash.CA2.p3[18] ;
 wire \hash.CA2.p3[19] ;
 wire \hash.CA2.p3[1] ;
 wire \hash.CA2.p3[20] ;
 wire \hash.CA2.p3[21] ;
 wire \hash.CA2.p3[22] ;
 wire \hash.CA2.p3[23] ;
 wire \hash.CA2.p3[24] ;
 wire \hash.CA2.p3[25] ;
 wire \hash.CA2.p3[26] ;
 wire \hash.CA2.p3[27] ;
 wire \hash.CA2.p3[28] ;
 wire \hash.CA2.p3[29] ;
 wire \hash.CA2.p3[2] ;
 wire \hash.CA2.p3[30] ;
 wire \hash.CA2.p3[31] ;
 wire \hash.CA2.p3[3] ;
 wire \hash.CA2.p3[4] ;
 wire \hash.CA2.p3[5] ;
 wire \hash.CA2.p3[6] ;
 wire \hash.CA2.p3[7] ;
 wire \hash.CA2.p3[8] ;
 wire \hash.CA2.p3[9] ;
 wire \hash.CA2.p4[0] ;
 wire \hash.CA2.p4[10] ;
 wire \hash.CA2.p4[11] ;
 wire \hash.CA2.p4[12] ;
 wire \hash.CA2.p4[13] ;
 wire \hash.CA2.p4[14] ;
 wire \hash.CA2.p4[15] ;
 wire \hash.CA2.p4[16] ;
 wire \hash.CA2.p4[17] ;
 wire \hash.CA2.p4[18] ;
 wire \hash.CA2.p4[19] ;
 wire \hash.CA2.p4[1] ;
 wire \hash.CA2.p4[20] ;
 wire \hash.CA2.p4[21] ;
 wire \hash.CA2.p4[22] ;
 wire \hash.CA2.p4[23] ;
 wire \hash.CA2.p4[24] ;
 wire \hash.CA2.p4[25] ;
 wire \hash.CA2.p4[26] ;
 wire \hash.CA2.p4[27] ;
 wire \hash.CA2.p4[28] ;
 wire \hash.CA2.p4[29] ;
 wire \hash.CA2.p4[2] ;
 wire \hash.CA2.p4[30] ;
 wire \hash.CA2.p4[31] ;
 wire \hash.CA2.p4[3] ;
 wire \hash.CA2.p4[4] ;
 wire \hash.CA2.p4[5] ;
 wire \hash.CA2.p4[6] ;
 wire \hash.CA2.p4[7] ;
 wire \hash.CA2.p4[8] ;
 wire \hash.CA2.p4[9] ;
 wire \hash.CA2.p5[0] ;
 wire \hash.CA2.p5[10] ;
 wire \hash.CA2.p5[11] ;
 wire \hash.CA2.p5[12] ;
 wire \hash.CA2.p5[13] ;
 wire \hash.CA2.p5[14] ;
 wire \hash.CA2.p5[15] ;
 wire \hash.CA2.p5[16] ;
 wire \hash.CA2.p5[17] ;
 wire \hash.CA2.p5[18] ;
 wire \hash.CA2.p5[19] ;
 wire \hash.CA2.p5[1] ;
 wire \hash.CA2.p5[20] ;
 wire \hash.CA2.p5[21] ;
 wire \hash.CA2.p5[22] ;
 wire \hash.CA2.p5[23] ;
 wire \hash.CA2.p5[24] ;
 wire \hash.CA2.p5[25] ;
 wire \hash.CA2.p5[26] ;
 wire \hash.CA2.p5[27] ;
 wire \hash.CA2.p5[28] ;
 wire \hash.CA2.p5[29] ;
 wire \hash.CA2.p5[2] ;
 wire \hash.CA2.p5[30] ;
 wire \hash.CA2.p5[31] ;
 wire \hash.CA2.p5[3] ;
 wire \hash.CA2.p5[4] ;
 wire \hash.CA2.p5[5] ;
 wire \hash.CA2.p5[6] ;
 wire \hash.CA2.p5[7] ;
 wire \hash.CA2.p5[8] ;
 wire \hash.CA2.p5[9] ;
 wire \hash.reset ;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire ready_dash;
 wire reset_hash;
 wire \w[0][0] ;
 wire \w[0][10] ;
 wire \w[0][11] ;
 wire \w[0][12] ;
 wire \w[0][13] ;
 wire \w[0][14] ;
 wire \w[0][15] ;
 wire \w[0][16] ;
 wire \w[0][17] ;
 wire \w[0][18] ;
 wire \w[0][19] ;
 wire \w[0][1] ;
 wire \w[0][20] ;
 wire \w[0][21] ;
 wire \w[0][22] ;
 wire \w[0][23] ;
 wire \w[0][24] ;
 wire \w[0][25] ;
 wire \w[0][26] ;
 wire \w[0][27] ;
 wire \w[0][28] ;
 wire \w[0][29] ;
 wire \w[0][2] ;
 wire \w[0][30] ;
 wire \w[0][31] ;
 wire \w[0][3] ;
 wire \w[0][4] ;
 wire \w[0][5] ;
 wire \w[0][6] ;
 wire \w[0][7] ;
 wire \w[0][8] ;
 wire \w[0][9] ;
 wire \w[10][0] ;
 wire \w[10][10] ;
 wire \w[10][11] ;
 wire \w[10][12] ;
 wire \w[10][13] ;
 wire \w[10][14] ;
 wire \w[10][15] ;
 wire \w[10][16] ;
 wire \w[10][17] ;
 wire \w[10][18] ;
 wire \w[10][19] ;
 wire \w[10][1] ;
 wire \w[10][20] ;
 wire \w[10][21] ;
 wire \w[10][22] ;
 wire \w[10][23] ;
 wire \w[10][24] ;
 wire \w[10][25] ;
 wire \w[10][26] ;
 wire \w[10][27] ;
 wire \w[10][28] ;
 wire \w[10][29] ;
 wire \w[10][2] ;
 wire \w[10][30] ;
 wire \w[10][31] ;
 wire \w[10][3] ;
 wire \w[10][4] ;
 wire \w[10][5] ;
 wire \w[10][6] ;
 wire \w[10][7] ;
 wire \w[10][8] ;
 wire \w[10][9] ;
 wire \w[11][0] ;
 wire \w[11][10] ;
 wire \w[11][11] ;
 wire \w[11][12] ;
 wire \w[11][13] ;
 wire \w[11][14] ;
 wire \w[11][15] ;
 wire \w[11][16] ;
 wire \w[11][17] ;
 wire \w[11][18] ;
 wire \w[11][19] ;
 wire \w[11][1] ;
 wire \w[11][20] ;
 wire \w[11][21] ;
 wire \w[11][22] ;
 wire \w[11][23] ;
 wire \w[11][24] ;
 wire \w[11][25] ;
 wire \w[11][26] ;
 wire \w[11][27] ;
 wire \w[11][28] ;
 wire \w[11][29] ;
 wire \w[11][2] ;
 wire \w[11][30] ;
 wire \w[11][31] ;
 wire \w[11][3] ;
 wire \w[11][4] ;
 wire \w[11][5] ;
 wire \w[11][6] ;
 wire \w[11][7] ;
 wire \w[11][8] ;
 wire \w[11][9] ;
 wire \w[12][0] ;
 wire \w[12][10] ;
 wire \w[12][11] ;
 wire \w[12][12] ;
 wire \w[12][13] ;
 wire \w[12][14] ;
 wire \w[12][15] ;
 wire \w[12][16] ;
 wire \w[12][17] ;
 wire \w[12][18] ;
 wire \w[12][19] ;
 wire \w[12][1] ;
 wire \w[12][20] ;
 wire \w[12][21] ;
 wire \w[12][22] ;
 wire \w[12][23] ;
 wire \w[12][24] ;
 wire \w[12][25] ;
 wire \w[12][26] ;
 wire \w[12][27] ;
 wire \w[12][28] ;
 wire \w[12][29] ;
 wire \w[12][2] ;
 wire \w[12][30] ;
 wire \w[12][31] ;
 wire \w[12][3] ;
 wire \w[12][4] ;
 wire \w[12][5] ;
 wire \w[12][6] ;
 wire \w[12][7] ;
 wire \w[12][8] ;
 wire \w[12][9] ;
 wire \w[13][0] ;
 wire \w[13][10] ;
 wire \w[13][11] ;
 wire \w[13][12] ;
 wire \w[13][13] ;
 wire \w[13][14] ;
 wire \w[13][15] ;
 wire \w[13][16] ;
 wire \w[13][17] ;
 wire \w[13][18] ;
 wire \w[13][19] ;
 wire \w[13][1] ;
 wire \w[13][20] ;
 wire \w[13][21] ;
 wire \w[13][22] ;
 wire \w[13][23] ;
 wire \w[13][24] ;
 wire \w[13][25] ;
 wire \w[13][26] ;
 wire \w[13][27] ;
 wire \w[13][28] ;
 wire \w[13][29] ;
 wire \w[13][2] ;
 wire \w[13][30] ;
 wire \w[13][31] ;
 wire \w[13][3] ;
 wire \w[13][4] ;
 wire \w[13][5] ;
 wire \w[13][6] ;
 wire \w[13][7] ;
 wire \w[13][8] ;
 wire \w[13][9] ;
 wire \w[14][0] ;
 wire \w[14][10] ;
 wire \w[14][11] ;
 wire \w[14][12] ;
 wire \w[14][13] ;
 wire \w[14][14] ;
 wire \w[14][15] ;
 wire \w[14][16] ;
 wire \w[14][17] ;
 wire \w[14][18] ;
 wire \w[14][19] ;
 wire \w[14][1] ;
 wire \w[14][20] ;
 wire \w[14][21] ;
 wire \w[14][22] ;
 wire \w[14][23] ;
 wire \w[14][24] ;
 wire \w[14][25] ;
 wire \w[14][26] ;
 wire \w[14][27] ;
 wire \w[14][28] ;
 wire \w[14][29] ;
 wire \w[14][2] ;
 wire \w[14][30] ;
 wire \w[14][31] ;
 wire \w[14][3] ;
 wire \w[14][4] ;
 wire \w[14][5] ;
 wire \w[14][6] ;
 wire \w[14][7] ;
 wire \w[14][8] ;
 wire \w[14][9] ;
 wire \w[15][0] ;
 wire \w[15][10] ;
 wire \w[15][11] ;
 wire \w[15][12] ;
 wire \w[15][13] ;
 wire \w[15][14] ;
 wire \w[15][15] ;
 wire \w[15][16] ;
 wire \w[15][17] ;
 wire \w[15][18] ;
 wire \w[15][19] ;
 wire \w[15][1] ;
 wire \w[15][20] ;
 wire \w[15][21] ;
 wire \w[15][22] ;
 wire \w[15][23] ;
 wire \w[15][24] ;
 wire \w[15][25] ;
 wire \w[15][26] ;
 wire \w[15][27] ;
 wire \w[15][28] ;
 wire \w[15][29] ;
 wire \w[15][2] ;
 wire \w[15][30] ;
 wire \w[15][31] ;
 wire \w[15][3] ;
 wire \w[15][4] ;
 wire \w[15][5] ;
 wire \w[15][6] ;
 wire \w[15][7] ;
 wire \w[15][8] ;
 wire \w[15][9] ;
 wire \w[16][0] ;
 wire \w[16][10] ;
 wire \w[16][11] ;
 wire \w[16][12] ;
 wire \w[16][13] ;
 wire \w[16][14] ;
 wire \w[16][15] ;
 wire \w[16][16] ;
 wire \w[16][17] ;
 wire \w[16][18] ;
 wire \w[16][19] ;
 wire \w[16][1] ;
 wire \w[16][20] ;
 wire \w[16][21] ;
 wire \w[16][22] ;
 wire \w[16][23] ;
 wire \w[16][24] ;
 wire \w[16][25] ;
 wire \w[16][26] ;
 wire \w[16][27] ;
 wire \w[16][28] ;
 wire \w[16][29] ;
 wire \w[16][2] ;
 wire \w[16][30] ;
 wire \w[16][31] ;
 wire \w[16][3] ;
 wire \w[16][4] ;
 wire \w[16][5] ;
 wire \w[16][6] ;
 wire \w[16][7] ;
 wire \w[16][8] ;
 wire \w[16][9] ;
 wire \w[17][0] ;
 wire \w[17][10] ;
 wire \w[17][11] ;
 wire \w[17][12] ;
 wire \w[17][13] ;
 wire \w[17][14] ;
 wire \w[17][15] ;
 wire \w[17][16] ;
 wire \w[17][17] ;
 wire \w[17][18] ;
 wire \w[17][19] ;
 wire \w[17][1] ;
 wire \w[17][20] ;
 wire \w[17][21] ;
 wire \w[17][22] ;
 wire \w[17][23] ;
 wire \w[17][24] ;
 wire \w[17][25] ;
 wire \w[17][26] ;
 wire \w[17][27] ;
 wire \w[17][28] ;
 wire \w[17][29] ;
 wire \w[17][2] ;
 wire \w[17][30] ;
 wire \w[17][31] ;
 wire \w[17][3] ;
 wire \w[17][4] ;
 wire \w[17][5] ;
 wire \w[17][6] ;
 wire \w[17][7] ;
 wire \w[17][8] ;
 wire \w[17][9] ;
 wire \w[18][0] ;
 wire \w[18][10] ;
 wire \w[18][11] ;
 wire \w[18][12] ;
 wire \w[18][13] ;
 wire \w[18][14] ;
 wire \w[18][15] ;
 wire \w[18][16] ;
 wire \w[18][17] ;
 wire \w[18][18] ;
 wire \w[18][19] ;
 wire \w[18][1] ;
 wire \w[18][20] ;
 wire \w[18][21] ;
 wire \w[18][22] ;
 wire \w[18][23] ;
 wire \w[18][24] ;
 wire \w[18][25] ;
 wire \w[18][26] ;
 wire \w[18][27] ;
 wire \w[18][28] ;
 wire \w[18][29] ;
 wire \w[18][2] ;
 wire \w[18][30] ;
 wire \w[18][31] ;
 wire \w[18][3] ;
 wire \w[18][4] ;
 wire \w[18][5] ;
 wire \w[18][6] ;
 wire \w[18][7] ;
 wire \w[18][8] ;
 wire \w[18][9] ;
 wire \w[19][0] ;
 wire \w[19][10] ;
 wire \w[19][11] ;
 wire \w[19][12] ;
 wire \w[19][13] ;
 wire \w[19][14] ;
 wire \w[19][15] ;
 wire \w[19][16] ;
 wire \w[19][17] ;
 wire \w[19][18] ;
 wire \w[19][19] ;
 wire \w[19][1] ;
 wire \w[19][20] ;
 wire \w[19][21] ;
 wire \w[19][22] ;
 wire \w[19][23] ;
 wire \w[19][24] ;
 wire \w[19][25] ;
 wire \w[19][26] ;
 wire \w[19][27] ;
 wire \w[19][28] ;
 wire \w[19][29] ;
 wire \w[19][2] ;
 wire \w[19][30] ;
 wire \w[19][31] ;
 wire \w[19][3] ;
 wire \w[19][4] ;
 wire \w[19][5] ;
 wire \w[19][6] ;
 wire \w[19][7] ;
 wire \w[19][8] ;
 wire \w[19][9] ;
 wire \w[1][0] ;
 wire \w[1][10] ;
 wire \w[1][11] ;
 wire \w[1][12] ;
 wire \w[1][13] ;
 wire \w[1][14] ;
 wire \w[1][15] ;
 wire \w[1][16] ;
 wire \w[1][17] ;
 wire \w[1][18] ;
 wire \w[1][19] ;
 wire \w[1][1] ;
 wire \w[1][20] ;
 wire \w[1][21] ;
 wire \w[1][22] ;
 wire \w[1][23] ;
 wire \w[1][24] ;
 wire \w[1][25] ;
 wire \w[1][26] ;
 wire \w[1][27] ;
 wire \w[1][28] ;
 wire \w[1][29] ;
 wire \w[1][2] ;
 wire \w[1][30] ;
 wire \w[1][31] ;
 wire \w[1][3] ;
 wire \w[1][4] ;
 wire \w[1][5] ;
 wire \w[1][6] ;
 wire \w[1][7] ;
 wire \w[1][8] ;
 wire \w[1][9] ;
 wire \w[20][0] ;
 wire \w[20][10] ;
 wire \w[20][11] ;
 wire \w[20][12] ;
 wire \w[20][13] ;
 wire \w[20][14] ;
 wire \w[20][15] ;
 wire \w[20][16] ;
 wire \w[20][17] ;
 wire \w[20][18] ;
 wire \w[20][19] ;
 wire \w[20][1] ;
 wire \w[20][20] ;
 wire \w[20][21] ;
 wire \w[20][22] ;
 wire \w[20][23] ;
 wire \w[20][24] ;
 wire \w[20][25] ;
 wire \w[20][26] ;
 wire \w[20][27] ;
 wire \w[20][28] ;
 wire \w[20][29] ;
 wire \w[20][2] ;
 wire \w[20][30] ;
 wire \w[20][31] ;
 wire \w[20][3] ;
 wire \w[20][4] ;
 wire \w[20][5] ;
 wire \w[20][6] ;
 wire \w[20][7] ;
 wire \w[20][8] ;
 wire \w[20][9] ;
 wire \w[21][0] ;
 wire \w[21][10] ;
 wire \w[21][11] ;
 wire \w[21][12] ;
 wire \w[21][13] ;
 wire \w[21][14] ;
 wire \w[21][15] ;
 wire \w[21][16] ;
 wire \w[21][17] ;
 wire \w[21][18] ;
 wire \w[21][19] ;
 wire \w[21][1] ;
 wire \w[21][20] ;
 wire \w[21][21] ;
 wire \w[21][22] ;
 wire \w[21][23] ;
 wire \w[21][24] ;
 wire \w[21][25] ;
 wire \w[21][26] ;
 wire \w[21][27] ;
 wire \w[21][28] ;
 wire \w[21][29] ;
 wire \w[21][2] ;
 wire \w[21][30] ;
 wire \w[21][31] ;
 wire \w[21][3] ;
 wire \w[21][4] ;
 wire \w[21][5] ;
 wire \w[21][6] ;
 wire \w[21][7] ;
 wire \w[21][8] ;
 wire \w[21][9] ;
 wire \w[22][0] ;
 wire \w[22][10] ;
 wire \w[22][11] ;
 wire \w[22][12] ;
 wire \w[22][13] ;
 wire \w[22][14] ;
 wire \w[22][15] ;
 wire \w[22][16] ;
 wire \w[22][17] ;
 wire \w[22][18] ;
 wire \w[22][19] ;
 wire \w[22][1] ;
 wire \w[22][20] ;
 wire \w[22][21] ;
 wire \w[22][22] ;
 wire \w[22][23] ;
 wire \w[22][24] ;
 wire \w[22][25] ;
 wire \w[22][26] ;
 wire \w[22][27] ;
 wire \w[22][28] ;
 wire \w[22][29] ;
 wire \w[22][2] ;
 wire \w[22][30] ;
 wire \w[22][31] ;
 wire \w[22][3] ;
 wire \w[22][4] ;
 wire \w[22][5] ;
 wire \w[22][6] ;
 wire \w[22][7] ;
 wire \w[22][8] ;
 wire \w[22][9] ;
 wire \w[23][0] ;
 wire \w[23][10] ;
 wire \w[23][11] ;
 wire \w[23][12] ;
 wire \w[23][13] ;
 wire \w[23][14] ;
 wire \w[23][15] ;
 wire \w[23][16] ;
 wire \w[23][17] ;
 wire \w[23][18] ;
 wire \w[23][19] ;
 wire \w[23][1] ;
 wire \w[23][20] ;
 wire \w[23][21] ;
 wire \w[23][22] ;
 wire \w[23][23] ;
 wire \w[23][24] ;
 wire \w[23][25] ;
 wire \w[23][26] ;
 wire \w[23][27] ;
 wire \w[23][28] ;
 wire \w[23][29] ;
 wire \w[23][2] ;
 wire \w[23][30] ;
 wire \w[23][31] ;
 wire \w[23][3] ;
 wire \w[23][4] ;
 wire \w[23][5] ;
 wire \w[23][6] ;
 wire \w[23][7] ;
 wire \w[23][8] ;
 wire \w[23][9] ;
 wire \w[24][0] ;
 wire \w[24][10] ;
 wire \w[24][11] ;
 wire \w[24][12] ;
 wire \w[24][13] ;
 wire \w[24][14] ;
 wire \w[24][15] ;
 wire \w[24][16] ;
 wire \w[24][17] ;
 wire \w[24][18] ;
 wire \w[24][19] ;
 wire \w[24][1] ;
 wire \w[24][20] ;
 wire \w[24][21] ;
 wire \w[24][22] ;
 wire \w[24][23] ;
 wire \w[24][24] ;
 wire \w[24][25] ;
 wire \w[24][26] ;
 wire \w[24][27] ;
 wire \w[24][28] ;
 wire \w[24][29] ;
 wire \w[24][2] ;
 wire \w[24][30] ;
 wire \w[24][31] ;
 wire \w[24][3] ;
 wire \w[24][4] ;
 wire \w[24][5] ;
 wire \w[24][6] ;
 wire \w[24][7] ;
 wire \w[24][8] ;
 wire \w[24][9] ;
 wire \w[25][0] ;
 wire \w[25][10] ;
 wire \w[25][11] ;
 wire \w[25][12] ;
 wire \w[25][13] ;
 wire \w[25][14] ;
 wire \w[25][15] ;
 wire \w[25][16] ;
 wire \w[25][17] ;
 wire \w[25][18] ;
 wire \w[25][19] ;
 wire \w[25][1] ;
 wire \w[25][20] ;
 wire \w[25][21] ;
 wire \w[25][22] ;
 wire \w[25][23] ;
 wire \w[25][24] ;
 wire \w[25][25] ;
 wire \w[25][26] ;
 wire \w[25][27] ;
 wire \w[25][28] ;
 wire \w[25][29] ;
 wire \w[25][2] ;
 wire \w[25][30] ;
 wire \w[25][31] ;
 wire \w[25][3] ;
 wire \w[25][4] ;
 wire \w[25][5] ;
 wire \w[25][6] ;
 wire \w[25][7] ;
 wire \w[25][8] ;
 wire \w[25][9] ;
 wire \w[26][0] ;
 wire \w[26][10] ;
 wire \w[26][11] ;
 wire \w[26][12] ;
 wire \w[26][13] ;
 wire \w[26][14] ;
 wire \w[26][15] ;
 wire \w[26][16] ;
 wire \w[26][17] ;
 wire \w[26][18] ;
 wire \w[26][19] ;
 wire \w[26][1] ;
 wire \w[26][20] ;
 wire \w[26][21] ;
 wire \w[26][22] ;
 wire \w[26][23] ;
 wire \w[26][24] ;
 wire \w[26][25] ;
 wire \w[26][26] ;
 wire \w[26][27] ;
 wire \w[26][28] ;
 wire \w[26][29] ;
 wire \w[26][2] ;
 wire \w[26][30] ;
 wire \w[26][31] ;
 wire \w[26][3] ;
 wire \w[26][4] ;
 wire \w[26][5] ;
 wire \w[26][6] ;
 wire \w[26][7] ;
 wire \w[26][8] ;
 wire \w[26][9] ;
 wire \w[27][0] ;
 wire \w[27][10] ;
 wire \w[27][11] ;
 wire \w[27][12] ;
 wire \w[27][13] ;
 wire \w[27][14] ;
 wire \w[27][15] ;
 wire \w[27][16] ;
 wire \w[27][17] ;
 wire \w[27][18] ;
 wire \w[27][19] ;
 wire \w[27][1] ;
 wire \w[27][20] ;
 wire \w[27][21] ;
 wire \w[27][22] ;
 wire \w[27][23] ;
 wire \w[27][24] ;
 wire \w[27][25] ;
 wire \w[27][26] ;
 wire \w[27][27] ;
 wire \w[27][28] ;
 wire \w[27][29] ;
 wire \w[27][2] ;
 wire \w[27][30] ;
 wire \w[27][31] ;
 wire \w[27][3] ;
 wire \w[27][4] ;
 wire \w[27][5] ;
 wire \w[27][6] ;
 wire \w[27][7] ;
 wire \w[27][8] ;
 wire \w[27][9] ;
 wire \w[28][0] ;
 wire \w[28][10] ;
 wire \w[28][11] ;
 wire \w[28][12] ;
 wire \w[28][13] ;
 wire \w[28][14] ;
 wire \w[28][15] ;
 wire \w[28][16] ;
 wire \w[28][17] ;
 wire \w[28][18] ;
 wire \w[28][19] ;
 wire \w[28][1] ;
 wire \w[28][20] ;
 wire \w[28][21] ;
 wire \w[28][22] ;
 wire \w[28][23] ;
 wire \w[28][24] ;
 wire \w[28][25] ;
 wire \w[28][26] ;
 wire \w[28][27] ;
 wire \w[28][28] ;
 wire \w[28][29] ;
 wire \w[28][2] ;
 wire \w[28][30] ;
 wire \w[28][31] ;
 wire \w[28][3] ;
 wire \w[28][4] ;
 wire \w[28][5] ;
 wire \w[28][6] ;
 wire \w[28][7] ;
 wire \w[28][8] ;
 wire \w[28][9] ;
 wire \w[29][0] ;
 wire \w[29][10] ;
 wire \w[29][11] ;
 wire \w[29][12] ;
 wire \w[29][13] ;
 wire \w[29][14] ;
 wire \w[29][15] ;
 wire \w[29][16] ;
 wire \w[29][17] ;
 wire \w[29][18] ;
 wire \w[29][19] ;
 wire \w[29][1] ;
 wire \w[29][20] ;
 wire \w[29][21] ;
 wire \w[29][22] ;
 wire \w[29][23] ;
 wire \w[29][24] ;
 wire \w[29][25] ;
 wire \w[29][26] ;
 wire \w[29][27] ;
 wire \w[29][28] ;
 wire \w[29][29] ;
 wire \w[29][2] ;
 wire \w[29][30] ;
 wire \w[29][31] ;
 wire \w[29][3] ;
 wire \w[29][4] ;
 wire \w[29][5] ;
 wire \w[29][6] ;
 wire \w[29][7] ;
 wire \w[29][8] ;
 wire \w[29][9] ;
 wire \w[2][0] ;
 wire \w[2][10] ;
 wire \w[2][11] ;
 wire \w[2][12] ;
 wire \w[2][13] ;
 wire \w[2][14] ;
 wire \w[2][15] ;
 wire \w[2][16] ;
 wire \w[2][17] ;
 wire \w[2][18] ;
 wire \w[2][19] ;
 wire \w[2][1] ;
 wire \w[2][20] ;
 wire \w[2][21] ;
 wire \w[2][22] ;
 wire \w[2][23] ;
 wire \w[2][24] ;
 wire \w[2][25] ;
 wire \w[2][26] ;
 wire \w[2][27] ;
 wire \w[2][28] ;
 wire \w[2][29] ;
 wire \w[2][2] ;
 wire \w[2][30] ;
 wire \w[2][31] ;
 wire \w[2][3] ;
 wire \w[2][4] ;
 wire \w[2][5] ;
 wire \w[2][6] ;
 wire \w[2][7] ;
 wire \w[2][8] ;
 wire \w[2][9] ;
 wire \w[30][0] ;
 wire \w[30][10] ;
 wire \w[30][11] ;
 wire \w[30][12] ;
 wire \w[30][13] ;
 wire \w[30][14] ;
 wire \w[30][15] ;
 wire \w[30][16] ;
 wire \w[30][17] ;
 wire \w[30][18] ;
 wire \w[30][19] ;
 wire \w[30][1] ;
 wire \w[30][20] ;
 wire \w[30][21] ;
 wire \w[30][22] ;
 wire \w[30][23] ;
 wire \w[30][24] ;
 wire \w[30][25] ;
 wire \w[30][26] ;
 wire \w[30][27] ;
 wire \w[30][28] ;
 wire \w[30][29] ;
 wire \w[30][2] ;
 wire \w[30][30] ;
 wire \w[30][31] ;
 wire \w[30][3] ;
 wire \w[30][4] ;
 wire \w[30][5] ;
 wire \w[30][6] ;
 wire \w[30][7] ;
 wire \w[30][8] ;
 wire \w[30][9] ;
 wire \w[31][0] ;
 wire \w[31][10] ;
 wire \w[31][11] ;
 wire \w[31][12] ;
 wire \w[31][13] ;
 wire \w[31][14] ;
 wire \w[31][15] ;
 wire \w[31][16] ;
 wire \w[31][17] ;
 wire \w[31][18] ;
 wire \w[31][19] ;
 wire \w[31][1] ;
 wire \w[31][20] ;
 wire \w[31][21] ;
 wire \w[31][22] ;
 wire \w[31][23] ;
 wire \w[31][24] ;
 wire \w[31][25] ;
 wire \w[31][26] ;
 wire \w[31][27] ;
 wire \w[31][28] ;
 wire \w[31][29] ;
 wire \w[31][2] ;
 wire \w[31][30] ;
 wire \w[31][31] ;
 wire \w[31][3] ;
 wire \w[31][4] ;
 wire \w[31][5] ;
 wire \w[31][6] ;
 wire \w[31][7] ;
 wire \w[31][8] ;
 wire \w[31][9] ;
 wire \w[32][0] ;
 wire \w[32][10] ;
 wire \w[32][11] ;
 wire \w[32][12] ;
 wire \w[32][13] ;
 wire \w[32][14] ;
 wire \w[32][15] ;
 wire \w[32][16] ;
 wire \w[32][17] ;
 wire \w[32][18] ;
 wire \w[32][19] ;
 wire \w[32][1] ;
 wire \w[32][20] ;
 wire \w[32][21] ;
 wire \w[32][22] ;
 wire \w[32][23] ;
 wire \w[32][24] ;
 wire \w[32][25] ;
 wire \w[32][26] ;
 wire \w[32][27] ;
 wire \w[32][28] ;
 wire \w[32][29] ;
 wire \w[32][2] ;
 wire \w[32][30] ;
 wire \w[32][31] ;
 wire \w[32][3] ;
 wire \w[32][4] ;
 wire \w[32][5] ;
 wire \w[32][6] ;
 wire \w[32][7] ;
 wire \w[32][8] ;
 wire \w[32][9] ;
 wire \w[33][0] ;
 wire \w[33][10] ;
 wire \w[33][11] ;
 wire \w[33][12] ;
 wire \w[33][13] ;
 wire \w[33][14] ;
 wire \w[33][15] ;
 wire \w[33][16] ;
 wire \w[33][17] ;
 wire \w[33][18] ;
 wire \w[33][19] ;
 wire \w[33][1] ;
 wire \w[33][20] ;
 wire \w[33][21] ;
 wire \w[33][22] ;
 wire \w[33][23] ;
 wire \w[33][24] ;
 wire \w[33][25] ;
 wire \w[33][26] ;
 wire \w[33][27] ;
 wire \w[33][28] ;
 wire \w[33][29] ;
 wire \w[33][2] ;
 wire \w[33][30] ;
 wire \w[33][31] ;
 wire \w[33][3] ;
 wire \w[33][4] ;
 wire \w[33][5] ;
 wire \w[33][6] ;
 wire \w[33][7] ;
 wire \w[33][8] ;
 wire \w[33][9] ;
 wire \w[34][0] ;
 wire \w[34][10] ;
 wire \w[34][11] ;
 wire \w[34][12] ;
 wire \w[34][13] ;
 wire \w[34][14] ;
 wire \w[34][15] ;
 wire \w[34][16] ;
 wire \w[34][17] ;
 wire \w[34][18] ;
 wire \w[34][19] ;
 wire \w[34][1] ;
 wire \w[34][20] ;
 wire \w[34][21] ;
 wire \w[34][22] ;
 wire \w[34][23] ;
 wire \w[34][24] ;
 wire \w[34][25] ;
 wire \w[34][26] ;
 wire \w[34][27] ;
 wire \w[34][28] ;
 wire \w[34][29] ;
 wire \w[34][2] ;
 wire \w[34][30] ;
 wire \w[34][31] ;
 wire \w[34][3] ;
 wire \w[34][4] ;
 wire \w[34][5] ;
 wire \w[34][6] ;
 wire \w[34][7] ;
 wire \w[34][8] ;
 wire \w[34][9] ;
 wire \w[35][0] ;
 wire \w[35][10] ;
 wire \w[35][11] ;
 wire \w[35][12] ;
 wire \w[35][13] ;
 wire \w[35][14] ;
 wire \w[35][15] ;
 wire \w[35][16] ;
 wire \w[35][17] ;
 wire \w[35][18] ;
 wire \w[35][19] ;
 wire \w[35][1] ;
 wire \w[35][20] ;
 wire \w[35][21] ;
 wire \w[35][22] ;
 wire \w[35][23] ;
 wire \w[35][24] ;
 wire \w[35][25] ;
 wire \w[35][26] ;
 wire \w[35][27] ;
 wire \w[35][28] ;
 wire \w[35][29] ;
 wire \w[35][2] ;
 wire \w[35][30] ;
 wire \w[35][31] ;
 wire \w[35][3] ;
 wire \w[35][4] ;
 wire \w[35][5] ;
 wire \w[35][6] ;
 wire \w[35][7] ;
 wire \w[35][8] ;
 wire \w[35][9] ;
 wire \w[36][0] ;
 wire \w[36][10] ;
 wire \w[36][11] ;
 wire \w[36][12] ;
 wire \w[36][13] ;
 wire \w[36][14] ;
 wire \w[36][15] ;
 wire \w[36][16] ;
 wire \w[36][17] ;
 wire \w[36][18] ;
 wire \w[36][19] ;
 wire \w[36][1] ;
 wire \w[36][20] ;
 wire \w[36][21] ;
 wire \w[36][22] ;
 wire \w[36][23] ;
 wire \w[36][24] ;
 wire \w[36][25] ;
 wire \w[36][26] ;
 wire \w[36][27] ;
 wire \w[36][28] ;
 wire \w[36][29] ;
 wire \w[36][2] ;
 wire \w[36][30] ;
 wire \w[36][31] ;
 wire \w[36][3] ;
 wire \w[36][4] ;
 wire \w[36][5] ;
 wire \w[36][6] ;
 wire \w[36][7] ;
 wire \w[36][8] ;
 wire \w[36][9] ;
 wire \w[37][0] ;
 wire \w[37][10] ;
 wire \w[37][11] ;
 wire \w[37][12] ;
 wire \w[37][13] ;
 wire \w[37][14] ;
 wire \w[37][15] ;
 wire \w[37][16] ;
 wire \w[37][17] ;
 wire \w[37][18] ;
 wire \w[37][19] ;
 wire \w[37][1] ;
 wire \w[37][20] ;
 wire \w[37][21] ;
 wire \w[37][22] ;
 wire \w[37][23] ;
 wire \w[37][24] ;
 wire \w[37][25] ;
 wire \w[37][26] ;
 wire \w[37][27] ;
 wire \w[37][28] ;
 wire \w[37][29] ;
 wire \w[37][2] ;
 wire \w[37][30] ;
 wire \w[37][31] ;
 wire \w[37][3] ;
 wire \w[37][4] ;
 wire \w[37][5] ;
 wire \w[37][6] ;
 wire \w[37][7] ;
 wire \w[37][8] ;
 wire \w[37][9] ;
 wire \w[38][0] ;
 wire \w[38][10] ;
 wire \w[38][11] ;
 wire \w[38][12] ;
 wire \w[38][13] ;
 wire \w[38][14] ;
 wire \w[38][15] ;
 wire \w[38][16] ;
 wire \w[38][17] ;
 wire \w[38][18] ;
 wire \w[38][19] ;
 wire \w[38][1] ;
 wire \w[38][20] ;
 wire \w[38][21] ;
 wire \w[38][22] ;
 wire \w[38][23] ;
 wire \w[38][24] ;
 wire \w[38][25] ;
 wire \w[38][26] ;
 wire \w[38][27] ;
 wire \w[38][28] ;
 wire \w[38][29] ;
 wire \w[38][2] ;
 wire \w[38][30] ;
 wire \w[38][31] ;
 wire \w[38][3] ;
 wire \w[38][4] ;
 wire \w[38][5] ;
 wire \w[38][6] ;
 wire \w[38][7] ;
 wire \w[38][8] ;
 wire \w[38][9] ;
 wire \w[39][0] ;
 wire \w[39][10] ;
 wire \w[39][11] ;
 wire \w[39][12] ;
 wire \w[39][13] ;
 wire \w[39][14] ;
 wire \w[39][15] ;
 wire \w[39][16] ;
 wire \w[39][17] ;
 wire \w[39][18] ;
 wire \w[39][19] ;
 wire \w[39][1] ;
 wire \w[39][20] ;
 wire \w[39][21] ;
 wire \w[39][22] ;
 wire \w[39][23] ;
 wire \w[39][24] ;
 wire \w[39][25] ;
 wire \w[39][26] ;
 wire \w[39][27] ;
 wire \w[39][28] ;
 wire \w[39][29] ;
 wire \w[39][2] ;
 wire \w[39][30] ;
 wire \w[39][31] ;
 wire \w[39][3] ;
 wire \w[39][4] ;
 wire \w[39][5] ;
 wire \w[39][6] ;
 wire \w[39][7] ;
 wire \w[39][8] ;
 wire \w[39][9] ;
 wire \w[3][0] ;
 wire \w[3][10] ;
 wire \w[3][11] ;
 wire \w[3][12] ;
 wire \w[3][13] ;
 wire \w[3][14] ;
 wire \w[3][15] ;
 wire \w[3][16] ;
 wire \w[3][17] ;
 wire \w[3][18] ;
 wire \w[3][19] ;
 wire \w[3][1] ;
 wire \w[3][20] ;
 wire \w[3][21] ;
 wire \w[3][22] ;
 wire \w[3][23] ;
 wire \w[3][24] ;
 wire \w[3][25] ;
 wire \w[3][26] ;
 wire \w[3][27] ;
 wire \w[3][28] ;
 wire \w[3][29] ;
 wire \w[3][2] ;
 wire \w[3][30] ;
 wire \w[3][31] ;
 wire \w[3][3] ;
 wire \w[3][4] ;
 wire \w[3][5] ;
 wire \w[3][6] ;
 wire \w[3][7] ;
 wire \w[3][8] ;
 wire \w[3][9] ;
 wire \w[40][0] ;
 wire \w[40][10] ;
 wire \w[40][11] ;
 wire \w[40][12] ;
 wire \w[40][13] ;
 wire \w[40][14] ;
 wire \w[40][15] ;
 wire \w[40][16] ;
 wire \w[40][17] ;
 wire \w[40][18] ;
 wire \w[40][19] ;
 wire \w[40][1] ;
 wire \w[40][20] ;
 wire \w[40][21] ;
 wire \w[40][22] ;
 wire \w[40][23] ;
 wire \w[40][24] ;
 wire \w[40][25] ;
 wire \w[40][26] ;
 wire \w[40][27] ;
 wire \w[40][28] ;
 wire \w[40][29] ;
 wire \w[40][2] ;
 wire \w[40][30] ;
 wire \w[40][31] ;
 wire \w[40][3] ;
 wire \w[40][4] ;
 wire \w[40][5] ;
 wire \w[40][6] ;
 wire \w[40][7] ;
 wire \w[40][8] ;
 wire \w[40][9] ;
 wire \w[41][0] ;
 wire \w[41][10] ;
 wire \w[41][11] ;
 wire \w[41][12] ;
 wire \w[41][13] ;
 wire \w[41][14] ;
 wire \w[41][15] ;
 wire \w[41][16] ;
 wire \w[41][17] ;
 wire \w[41][18] ;
 wire \w[41][19] ;
 wire \w[41][1] ;
 wire \w[41][20] ;
 wire \w[41][21] ;
 wire \w[41][22] ;
 wire \w[41][23] ;
 wire \w[41][24] ;
 wire \w[41][25] ;
 wire \w[41][26] ;
 wire \w[41][27] ;
 wire \w[41][28] ;
 wire \w[41][29] ;
 wire \w[41][2] ;
 wire \w[41][30] ;
 wire \w[41][31] ;
 wire \w[41][3] ;
 wire \w[41][4] ;
 wire \w[41][5] ;
 wire \w[41][6] ;
 wire \w[41][7] ;
 wire \w[41][8] ;
 wire \w[41][9] ;
 wire \w[42][0] ;
 wire \w[42][10] ;
 wire \w[42][11] ;
 wire \w[42][12] ;
 wire \w[42][13] ;
 wire \w[42][14] ;
 wire \w[42][15] ;
 wire \w[42][16] ;
 wire \w[42][17] ;
 wire \w[42][18] ;
 wire \w[42][19] ;
 wire \w[42][1] ;
 wire \w[42][20] ;
 wire \w[42][21] ;
 wire \w[42][22] ;
 wire \w[42][23] ;
 wire \w[42][24] ;
 wire \w[42][25] ;
 wire \w[42][26] ;
 wire \w[42][27] ;
 wire \w[42][28] ;
 wire \w[42][29] ;
 wire \w[42][2] ;
 wire \w[42][30] ;
 wire \w[42][31] ;
 wire \w[42][3] ;
 wire \w[42][4] ;
 wire \w[42][5] ;
 wire \w[42][6] ;
 wire \w[42][7] ;
 wire \w[42][8] ;
 wire \w[42][9] ;
 wire \w[43][0] ;
 wire \w[43][10] ;
 wire \w[43][11] ;
 wire \w[43][12] ;
 wire \w[43][13] ;
 wire \w[43][14] ;
 wire \w[43][15] ;
 wire \w[43][16] ;
 wire \w[43][17] ;
 wire \w[43][18] ;
 wire \w[43][19] ;
 wire \w[43][1] ;
 wire \w[43][20] ;
 wire \w[43][21] ;
 wire \w[43][22] ;
 wire \w[43][23] ;
 wire \w[43][24] ;
 wire \w[43][25] ;
 wire \w[43][26] ;
 wire \w[43][27] ;
 wire \w[43][28] ;
 wire \w[43][29] ;
 wire \w[43][2] ;
 wire \w[43][30] ;
 wire \w[43][31] ;
 wire \w[43][3] ;
 wire \w[43][4] ;
 wire \w[43][5] ;
 wire \w[43][6] ;
 wire \w[43][7] ;
 wire \w[43][8] ;
 wire \w[43][9] ;
 wire \w[44][0] ;
 wire \w[44][10] ;
 wire \w[44][11] ;
 wire \w[44][12] ;
 wire \w[44][13] ;
 wire \w[44][14] ;
 wire \w[44][15] ;
 wire \w[44][16] ;
 wire \w[44][17] ;
 wire \w[44][18] ;
 wire \w[44][19] ;
 wire \w[44][1] ;
 wire \w[44][20] ;
 wire \w[44][21] ;
 wire \w[44][22] ;
 wire \w[44][23] ;
 wire \w[44][24] ;
 wire \w[44][25] ;
 wire \w[44][26] ;
 wire \w[44][27] ;
 wire \w[44][28] ;
 wire \w[44][29] ;
 wire \w[44][2] ;
 wire \w[44][30] ;
 wire \w[44][31] ;
 wire \w[44][3] ;
 wire \w[44][4] ;
 wire \w[44][5] ;
 wire \w[44][6] ;
 wire \w[44][7] ;
 wire \w[44][8] ;
 wire \w[44][9] ;
 wire \w[45][0] ;
 wire \w[45][10] ;
 wire \w[45][11] ;
 wire \w[45][12] ;
 wire \w[45][13] ;
 wire \w[45][14] ;
 wire \w[45][15] ;
 wire \w[45][16] ;
 wire \w[45][17] ;
 wire \w[45][18] ;
 wire \w[45][19] ;
 wire \w[45][1] ;
 wire \w[45][20] ;
 wire \w[45][21] ;
 wire \w[45][22] ;
 wire \w[45][23] ;
 wire \w[45][24] ;
 wire \w[45][25] ;
 wire \w[45][26] ;
 wire \w[45][27] ;
 wire \w[45][28] ;
 wire \w[45][29] ;
 wire \w[45][2] ;
 wire \w[45][30] ;
 wire \w[45][31] ;
 wire \w[45][3] ;
 wire \w[45][4] ;
 wire \w[45][5] ;
 wire \w[45][6] ;
 wire \w[45][7] ;
 wire \w[45][8] ;
 wire \w[45][9] ;
 wire \w[46][0] ;
 wire \w[46][10] ;
 wire \w[46][11] ;
 wire \w[46][12] ;
 wire \w[46][13] ;
 wire \w[46][14] ;
 wire \w[46][15] ;
 wire \w[46][16] ;
 wire \w[46][17] ;
 wire \w[46][18] ;
 wire \w[46][19] ;
 wire \w[46][1] ;
 wire \w[46][20] ;
 wire \w[46][21] ;
 wire \w[46][22] ;
 wire \w[46][23] ;
 wire \w[46][24] ;
 wire \w[46][25] ;
 wire \w[46][26] ;
 wire \w[46][27] ;
 wire \w[46][28] ;
 wire \w[46][29] ;
 wire \w[46][2] ;
 wire \w[46][30] ;
 wire \w[46][31] ;
 wire \w[46][3] ;
 wire \w[46][4] ;
 wire \w[46][5] ;
 wire \w[46][6] ;
 wire \w[46][7] ;
 wire \w[46][8] ;
 wire \w[46][9] ;
 wire \w[47][0] ;
 wire \w[47][10] ;
 wire \w[47][11] ;
 wire \w[47][12] ;
 wire \w[47][13] ;
 wire \w[47][14] ;
 wire \w[47][15] ;
 wire \w[47][16] ;
 wire \w[47][17] ;
 wire \w[47][18] ;
 wire \w[47][19] ;
 wire \w[47][1] ;
 wire \w[47][20] ;
 wire \w[47][21] ;
 wire \w[47][22] ;
 wire \w[47][23] ;
 wire \w[47][24] ;
 wire \w[47][25] ;
 wire \w[47][26] ;
 wire \w[47][27] ;
 wire \w[47][28] ;
 wire \w[47][29] ;
 wire \w[47][2] ;
 wire \w[47][30] ;
 wire \w[47][31] ;
 wire \w[47][3] ;
 wire \w[47][4] ;
 wire \w[47][5] ;
 wire \w[47][6] ;
 wire \w[47][7] ;
 wire \w[47][8] ;
 wire \w[47][9] ;
 wire \w[48][0] ;
 wire \w[48][10] ;
 wire \w[48][11] ;
 wire \w[48][12] ;
 wire \w[48][13] ;
 wire \w[48][14] ;
 wire \w[48][15] ;
 wire \w[48][16] ;
 wire \w[48][17] ;
 wire \w[48][18] ;
 wire \w[48][19] ;
 wire \w[48][1] ;
 wire \w[48][20] ;
 wire \w[48][21] ;
 wire \w[48][22] ;
 wire \w[48][23] ;
 wire \w[48][24] ;
 wire \w[48][25] ;
 wire \w[48][26] ;
 wire \w[48][27] ;
 wire \w[48][28] ;
 wire \w[48][29] ;
 wire \w[48][2] ;
 wire \w[48][30] ;
 wire \w[48][31] ;
 wire \w[48][3] ;
 wire \w[48][4] ;
 wire \w[48][5] ;
 wire \w[48][6] ;
 wire \w[48][7] ;
 wire \w[48][8] ;
 wire \w[48][9] ;
 wire \w[49][0] ;
 wire \w[49][10] ;
 wire \w[49][11] ;
 wire \w[49][12] ;
 wire \w[49][13] ;
 wire \w[49][14] ;
 wire \w[49][15] ;
 wire \w[49][16] ;
 wire \w[49][17] ;
 wire \w[49][18] ;
 wire \w[49][19] ;
 wire \w[49][1] ;
 wire \w[49][20] ;
 wire \w[49][21] ;
 wire \w[49][22] ;
 wire \w[49][23] ;
 wire \w[49][24] ;
 wire \w[49][25] ;
 wire \w[49][26] ;
 wire \w[49][27] ;
 wire \w[49][28] ;
 wire \w[49][29] ;
 wire \w[49][2] ;
 wire \w[49][30] ;
 wire \w[49][31] ;
 wire \w[49][3] ;
 wire \w[49][4] ;
 wire \w[49][5] ;
 wire \w[49][6] ;
 wire \w[49][7] ;
 wire \w[49][8] ;
 wire \w[49][9] ;
 wire \w[4][0] ;
 wire \w[4][10] ;
 wire \w[4][11] ;
 wire \w[4][12] ;
 wire \w[4][13] ;
 wire \w[4][14] ;
 wire \w[4][15] ;
 wire \w[4][16] ;
 wire \w[4][17] ;
 wire \w[4][18] ;
 wire \w[4][19] ;
 wire \w[4][1] ;
 wire \w[4][20] ;
 wire \w[4][21] ;
 wire \w[4][22] ;
 wire \w[4][23] ;
 wire \w[4][24] ;
 wire \w[4][25] ;
 wire \w[4][26] ;
 wire \w[4][27] ;
 wire \w[4][28] ;
 wire \w[4][29] ;
 wire \w[4][2] ;
 wire \w[4][30] ;
 wire \w[4][31] ;
 wire \w[4][3] ;
 wire \w[4][4] ;
 wire \w[4][5] ;
 wire \w[4][6] ;
 wire \w[4][7] ;
 wire \w[4][8] ;
 wire \w[4][9] ;
 wire \w[50][0] ;
 wire \w[50][10] ;
 wire \w[50][11] ;
 wire \w[50][12] ;
 wire \w[50][13] ;
 wire \w[50][14] ;
 wire \w[50][15] ;
 wire \w[50][16] ;
 wire \w[50][17] ;
 wire \w[50][18] ;
 wire \w[50][19] ;
 wire \w[50][1] ;
 wire \w[50][20] ;
 wire \w[50][21] ;
 wire \w[50][22] ;
 wire \w[50][23] ;
 wire \w[50][24] ;
 wire \w[50][25] ;
 wire \w[50][26] ;
 wire \w[50][27] ;
 wire \w[50][28] ;
 wire \w[50][29] ;
 wire \w[50][2] ;
 wire \w[50][30] ;
 wire \w[50][31] ;
 wire \w[50][3] ;
 wire \w[50][4] ;
 wire \w[50][5] ;
 wire \w[50][6] ;
 wire \w[50][7] ;
 wire \w[50][8] ;
 wire \w[50][9] ;
 wire \w[51][0] ;
 wire \w[51][10] ;
 wire \w[51][11] ;
 wire \w[51][12] ;
 wire \w[51][13] ;
 wire \w[51][14] ;
 wire \w[51][15] ;
 wire \w[51][16] ;
 wire \w[51][17] ;
 wire \w[51][18] ;
 wire \w[51][19] ;
 wire \w[51][1] ;
 wire \w[51][20] ;
 wire \w[51][21] ;
 wire \w[51][22] ;
 wire \w[51][23] ;
 wire \w[51][24] ;
 wire \w[51][25] ;
 wire \w[51][26] ;
 wire \w[51][27] ;
 wire \w[51][28] ;
 wire \w[51][29] ;
 wire \w[51][2] ;
 wire \w[51][30] ;
 wire \w[51][31] ;
 wire \w[51][3] ;
 wire \w[51][4] ;
 wire \w[51][5] ;
 wire \w[51][6] ;
 wire \w[51][7] ;
 wire \w[51][8] ;
 wire \w[51][9] ;
 wire \w[52][0] ;
 wire \w[52][10] ;
 wire \w[52][11] ;
 wire \w[52][12] ;
 wire \w[52][13] ;
 wire \w[52][14] ;
 wire \w[52][15] ;
 wire \w[52][16] ;
 wire \w[52][17] ;
 wire \w[52][18] ;
 wire \w[52][19] ;
 wire \w[52][1] ;
 wire \w[52][20] ;
 wire \w[52][21] ;
 wire \w[52][22] ;
 wire \w[52][23] ;
 wire \w[52][24] ;
 wire \w[52][25] ;
 wire \w[52][26] ;
 wire \w[52][27] ;
 wire \w[52][28] ;
 wire \w[52][29] ;
 wire \w[52][2] ;
 wire \w[52][30] ;
 wire \w[52][31] ;
 wire \w[52][3] ;
 wire \w[52][4] ;
 wire \w[52][5] ;
 wire \w[52][6] ;
 wire \w[52][7] ;
 wire \w[52][8] ;
 wire \w[52][9] ;
 wire \w[53][0] ;
 wire \w[53][10] ;
 wire \w[53][11] ;
 wire \w[53][12] ;
 wire \w[53][13] ;
 wire \w[53][14] ;
 wire \w[53][15] ;
 wire \w[53][16] ;
 wire \w[53][17] ;
 wire \w[53][18] ;
 wire \w[53][19] ;
 wire \w[53][1] ;
 wire \w[53][20] ;
 wire \w[53][21] ;
 wire \w[53][22] ;
 wire \w[53][23] ;
 wire \w[53][24] ;
 wire \w[53][25] ;
 wire \w[53][26] ;
 wire \w[53][27] ;
 wire \w[53][28] ;
 wire \w[53][29] ;
 wire \w[53][2] ;
 wire \w[53][30] ;
 wire \w[53][31] ;
 wire \w[53][3] ;
 wire \w[53][4] ;
 wire \w[53][5] ;
 wire \w[53][6] ;
 wire \w[53][7] ;
 wire \w[53][8] ;
 wire \w[53][9] ;
 wire \w[54][0] ;
 wire \w[54][10] ;
 wire \w[54][11] ;
 wire \w[54][12] ;
 wire \w[54][13] ;
 wire \w[54][14] ;
 wire \w[54][15] ;
 wire \w[54][16] ;
 wire \w[54][17] ;
 wire \w[54][18] ;
 wire \w[54][19] ;
 wire \w[54][1] ;
 wire \w[54][20] ;
 wire \w[54][21] ;
 wire \w[54][22] ;
 wire \w[54][23] ;
 wire \w[54][24] ;
 wire \w[54][25] ;
 wire \w[54][26] ;
 wire \w[54][27] ;
 wire \w[54][28] ;
 wire \w[54][29] ;
 wire \w[54][2] ;
 wire \w[54][30] ;
 wire \w[54][31] ;
 wire \w[54][3] ;
 wire \w[54][4] ;
 wire \w[54][5] ;
 wire \w[54][6] ;
 wire \w[54][7] ;
 wire \w[54][8] ;
 wire \w[54][9] ;
 wire \w[55][0] ;
 wire \w[55][10] ;
 wire \w[55][11] ;
 wire \w[55][12] ;
 wire \w[55][13] ;
 wire \w[55][14] ;
 wire \w[55][15] ;
 wire \w[55][16] ;
 wire \w[55][17] ;
 wire \w[55][18] ;
 wire \w[55][19] ;
 wire \w[55][1] ;
 wire \w[55][20] ;
 wire \w[55][21] ;
 wire \w[55][22] ;
 wire \w[55][23] ;
 wire \w[55][24] ;
 wire \w[55][25] ;
 wire \w[55][26] ;
 wire \w[55][27] ;
 wire \w[55][28] ;
 wire \w[55][29] ;
 wire \w[55][2] ;
 wire \w[55][30] ;
 wire \w[55][31] ;
 wire \w[55][3] ;
 wire \w[55][4] ;
 wire \w[55][5] ;
 wire \w[55][6] ;
 wire \w[55][7] ;
 wire \w[55][8] ;
 wire \w[55][9] ;
 wire \w[56][0] ;
 wire \w[56][10] ;
 wire \w[56][11] ;
 wire \w[56][12] ;
 wire \w[56][13] ;
 wire \w[56][14] ;
 wire \w[56][15] ;
 wire \w[56][16] ;
 wire \w[56][17] ;
 wire \w[56][18] ;
 wire \w[56][19] ;
 wire \w[56][1] ;
 wire \w[56][20] ;
 wire \w[56][21] ;
 wire \w[56][22] ;
 wire \w[56][23] ;
 wire \w[56][24] ;
 wire \w[56][25] ;
 wire \w[56][26] ;
 wire \w[56][27] ;
 wire \w[56][28] ;
 wire \w[56][29] ;
 wire \w[56][2] ;
 wire \w[56][30] ;
 wire \w[56][31] ;
 wire \w[56][3] ;
 wire \w[56][4] ;
 wire \w[56][5] ;
 wire \w[56][6] ;
 wire \w[56][7] ;
 wire \w[56][8] ;
 wire \w[56][9] ;
 wire \w[57][0] ;
 wire \w[57][10] ;
 wire \w[57][11] ;
 wire \w[57][12] ;
 wire \w[57][13] ;
 wire \w[57][14] ;
 wire \w[57][15] ;
 wire \w[57][16] ;
 wire \w[57][17] ;
 wire \w[57][18] ;
 wire \w[57][19] ;
 wire \w[57][1] ;
 wire \w[57][20] ;
 wire \w[57][21] ;
 wire \w[57][22] ;
 wire \w[57][23] ;
 wire \w[57][24] ;
 wire \w[57][25] ;
 wire \w[57][26] ;
 wire \w[57][27] ;
 wire \w[57][28] ;
 wire \w[57][29] ;
 wire \w[57][2] ;
 wire \w[57][30] ;
 wire \w[57][31] ;
 wire \w[57][3] ;
 wire \w[57][4] ;
 wire \w[57][5] ;
 wire \w[57][6] ;
 wire \w[57][7] ;
 wire \w[57][8] ;
 wire \w[57][9] ;
 wire \w[58][0] ;
 wire \w[58][10] ;
 wire \w[58][11] ;
 wire \w[58][12] ;
 wire \w[58][13] ;
 wire \w[58][14] ;
 wire \w[58][15] ;
 wire \w[58][16] ;
 wire \w[58][17] ;
 wire \w[58][18] ;
 wire \w[58][19] ;
 wire \w[58][1] ;
 wire \w[58][20] ;
 wire \w[58][21] ;
 wire \w[58][22] ;
 wire \w[58][23] ;
 wire \w[58][24] ;
 wire \w[58][25] ;
 wire \w[58][26] ;
 wire \w[58][27] ;
 wire \w[58][28] ;
 wire \w[58][29] ;
 wire \w[58][2] ;
 wire \w[58][30] ;
 wire \w[58][31] ;
 wire \w[58][3] ;
 wire \w[58][4] ;
 wire \w[58][5] ;
 wire \w[58][6] ;
 wire \w[58][7] ;
 wire \w[58][8] ;
 wire \w[58][9] ;
 wire \w[59][0] ;
 wire \w[59][10] ;
 wire \w[59][11] ;
 wire \w[59][12] ;
 wire \w[59][13] ;
 wire \w[59][14] ;
 wire \w[59][15] ;
 wire \w[59][16] ;
 wire \w[59][17] ;
 wire \w[59][18] ;
 wire \w[59][19] ;
 wire \w[59][1] ;
 wire \w[59][20] ;
 wire \w[59][21] ;
 wire \w[59][22] ;
 wire \w[59][23] ;
 wire \w[59][24] ;
 wire \w[59][25] ;
 wire \w[59][26] ;
 wire \w[59][27] ;
 wire \w[59][28] ;
 wire \w[59][29] ;
 wire \w[59][2] ;
 wire \w[59][30] ;
 wire \w[59][31] ;
 wire \w[59][3] ;
 wire \w[59][4] ;
 wire \w[59][5] ;
 wire \w[59][6] ;
 wire \w[59][7] ;
 wire \w[59][8] ;
 wire \w[59][9] ;
 wire \w[5][0] ;
 wire \w[5][10] ;
 wire \w[5][11] ;
 wire \w[5][12] ;
 wire \w[5][13] ;
 wire \w[5][14] ;
 wire \w[5][15] ;
 wire \w[5][16] ;
 wire \w[5][17] ;
 wire \w[5][18] ;
 wire \w[5][19] ;
 wire \w[5][1] ;
 wire \w[5][20] ;
 wire \w[5][21] ;
 wire \w[5][22] ;
 wire \w[5][23] ;
 wire \w[5][24] ;
 wire \w[5][25] ;
 wire \w[5][26] ;
 wire \w[5][27] ;
 wire \w[5][28] ;
 wire \w[5][29] ;
 wire \w[5][2] ;
 wire \w[5][30] ;
 wire \w[5][31] ;
 wire \w[5][3] ;
 wire \w[5][4] ;
 wire \w[5][5] ;
 wire \w[5][6] ;
 wire \w[5][7] ;
 wire \w[5][8] ;
 wire \w[5][9] ;
 wire \w[60][0] ;
 wire \w[60][10] ;
 wire \w[60][11] ;
 wire \w[60][12] ;
 wire \w[60][13] ;
 wire \w[60][14] ;
 wire \w[60][15] ;
 wire \w[60][16] ;
 wire \w[60][17] ;
 wire \w[60][18] ;
 wire \w[60][19] ;
 wire \w[60][1] ;
 wire \w[60][20] ;
 wire \w[60][21] ;
 wire \w[60][22] ;
 wire \w[60][23] ;
 wire \w[60][24] ;
 wire \w[60][25] ;
 wire \w[60][26] ;
 wire \w[60][27] ;
 wire \w[60][28] ;
 wire \w[60][29] ;
 wire \w[60][2] ;
 wire \w[60][30] ;
 wire \w[60][31] ;
 wire \w[60][3] ;
 wire \w[60][4] ;
 wire \w[60][5] ;
 wire \w[60][6] ;
 wire \w[60][7] ;
 wire \w[60][8] ;
 wire \w[60][9] ;
 wire \w[61][0] ;
 wire \w[61][10] ;
 wire \w[61][11] ;
 wire \w[61][12] ;
 wire \w[61][13] ;
 wire \w[61][14] ;
 wire \w[61][15] ;
 wire \w[61][16] ;
 wire \w[61][17] ;
 wire \w[61][18] ;
 wire \w[61][19] ;
 wire \w[61][1] ;
 wire \w[61][20] ;
 wire \w[61][21] ;
 wire \w[61][22] ;
 wire \w[61][23] ;
 wire \w[61][24] ;
 wire \w[61][25] ;
 wire \w[61][26] ;
 wire \w[61][27] ;
 wire \w[61][28] ;
 wire \w[61][29] ;
 wire \w[61][2] ;
 wire \w[61][30] ;
 wire \w[61][31] ;
 wire \w[61][3] ;
 wire \w[61][4] ;
 wire \w[61][5] ;
 wire \w[61][6] ;
 wire \w[61][7] ;
 wire \w[61][8] ;
 wire \w[61][9] ;
 wire \w[62][0] ;
 wire \w[62][10] ;
 wire \w[62][11] ;
 wire \w[62][12] ;
 wire \w[62][13] ;
 wire \w[62][14] ;
 wire \w[62][15] ;
 wire \w[62][16] ;
 wire \w[62][17] ;
 wire \w[62][18] ;
 wire \w[62][19] ;
 wire \w[62][1] ;
 wire \w[62][20] ;
 wire \w[62][21] ;
 wire \w[62][22] ;
 wire \w[62][23] ;
 wire \w[62][24] ;
 wire \w[62][25] ;
 wire \w[62][26] ;
 wire \w[62][27] ;
 wire \w[62][28] ;
 wire \w[62][29] ;
 wire \w[62][2] ;
 wire \w[62][30] ;
 wire \w[62][31] ;
 wire \w[62][3] ;
 wire \w[62][4] ;
 wire \w[62][5] ;
 wire \w[62][6] ;
 wire \w[62][7] ;
 wire \w[62][8] ;
 wire \w[62][9] ;
 wire \w[63][0] ;
 wire \w[63][10] ;
 wire \w[63][11] ;
 wire \w[63][12] ;
 wire \w[63][13] ;
 wire \w[63][14] ;
 wire \w[63][15] ;
 wire \w[63][16] ;
 wire \w[63][17] ;
 wire \w[63][18] ;
 wire \w[63][19] ;
 wire \w[63][1] ;
 wire \w[63][20] ;
 wire \w[63][21] ;
 wire \w[63][22] ;
 wire \w[63][23] ;
 wire \w[63][24] ;
 wire \w[63][25] ;
 wire \w[63][26] ;
 wire \w[63][27] ;
 wire \w[63][28] ;
 wire \w[63][29] ;
 wire \w[63][2] ;
 wire \w[63][30] ;
 wire \w[63][31] ;
 wire \w[63][3] ;
 wire \w[63][4] ;
 wire \w[63][5] ;
 wire \w[63][6] ;
 wire \w[63][7] ;
 wire \w[63][8] ;
 wire \w[63][9] ;
 wire \w[6][0] ;
 wire \w[6][10] ;
 wire \w[6][11] ;
 wire \w[6][12] ;
 wire \w[6][13] ;
 wire \w[6][14] ;
 wire \w[6][15] ;
 wire \w[6][16] ;
 wire \w[6][17] ;
 wire \w[6][18] ;
 wire \w[6][19] ;
 wire \w[6][1] ;
 wire \w[6][20] ;
 wire \w[6][21] ;
 wire \w[6][22] ;
 wire \w[6][23] ;
 wire \w[6][24] ;
 wire \w[6][25] ;
 wire \w[6][26] ;
 wire \w[6][27] ;
 wire \w[6][28] ;
 wire \w[6][29] ;
 wire \w[6][2] ;
 wire \w[6][30] ;
 wire \w[6][31] ;
 wire \w[6][3] ;
 wire \w[6][4] ;
 wire \w[6][5] ;
 wire \w[6][6] ;
 wire \w[6][7] ;
 wire \w[6][8] ;
 wire \w[6][9] ;
 wire \w[7][0] ;
 wire \w[7][10] ;
 wire \w[7][11] ;
 wire \w[7][12] ;
 wire \w[7][13] ;
 wire \w[7][14] ;
 wire \w[7][15] ;
 wire \w[7][16] ;
 wire \w[7][17] ;
 wire \w[7][18] ;
 wire \w[7][19] ;
 wire \w[7][1] ;
 wire \w[7][20] ;
 wire \w[7][21] ;
 wire \w[7][22] ;
 wire \w[7][23] ;
 wire \w[7][24] ;
 wire \w[7][25] ;
 wire \w[7][26] ;
 wire \w[7][27] ;
 wire \w[7][28] ;
 wire \w[7][29] ;
 wire \w[7][2] ;
 wire \w[7][30] ;
 wire \w[7][31] ;
 wire \w[7][3] ;
 wire \w[7][4] ;
 wire \w[7][5] ;
 wire \w[7][6] ;
 wire \w[7][7] ;
 wire \w[7][8] ;
 wire \w[7][9] ;
 wire \w[8][0] ;
 wire \w[8][10] ;
 wire \w[8][11] ;
 wire \w[8][12] ;
 wire \w[8][13] ;
 wire \w[8][14] ;
 wire \w[8][15] ;
 wire \w[8][16] ;
 wire \w[8][17] ;
 wire \w[8][18] ;
 wire \w[8][19] ;
 wire \w[8][1] ;
 wire \w[8][20] ;
 wire \w[8][21] ;
 wire \w[8][22] ;
 wire \w[8][23] ;
 wire \w[8][24] ;
 wire \w[8][25] ;
 wire \w[8][26] ;
 wire \w[8][27] ;
 wire \w[8][28] ;
 wire \w[8][29] ;
 wire \w[8][2] ;
 wire \w[8][30] ;
 wire \w[8][31] ;
 wire \w[8][3] ;
 wire \w[8][4] ;
 wire \w[8][5] ;
 wire \w[8][6] ;
 wire \w[8][7] ;
 wire \w[8][8] ;
 wire \w[8][9] ;
 wire \w[9][0] ;
 wire \w[9][10] ;
 wire \w[9][11] ;
 wire \w[9][12] ;
 wire \w[9][13] ;
 wire \w[9][14] ;
 wire \w[9][15] ;
 wire \w[9][16] ;
 wire \w[9][17] ;
 wire \w[9][18] ;
 wire \w[9][19] ;
 wire \w[9][1] ;
 wire \w[9][20] ;
 wire \w[9][21] ;
 wire \w[9][22] ;
 wire \w[9][23] ;
 wire \w[9][24] ;
 wire \w[9][25] ;
 wire \w[9][26] ;
 wire \w[9][27] ;
 wire \w[9][28] ;
 wire \w[9][29] ;
 wire \w[9][2] ;
 wire \w[9][30] ;
 wire \w[9][31] ;
 wire \w[9][3] ;
 wire \w[9][4] ;
 wire \w[9][5] ;
 wire \w[9][6] ;
 wire \w[9][7] ;
 wire \w[9][8] ;
 wire \w[9][9] ;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;

 sky130_fd_sc_hd__mux4_2 _14209_ (.A0(\w[33][14] ),
    .A1(\w[37][14] ),
    .A2(\w[35][14] ),
    .A3(\w[39][14] ),
    .S0(net465),
    .S1(net468),
    .X(_03883_));
 sky130_fd_sc_hd__mux4_2 _14210_ (.A0(\w[41][14] ),
    .A1(\w[45][14] ),
    .A2(\w[43][14] ),
    .A3(\w[47][14] ),
    .S0(net465),
    .S1(net468),
    .X(_03884_));
 sky130_fd_sc_hd__mux4_2 _14211_ (.A0(\w[49][14] ),
    .A1(\w[53][14] ),
    .A2(\w[51][14] ),
    .A3(\w[55][14] ),
    .S0(net465),
    .S1(net468),
    .X(_03885_));
 sky130_fd_sc_hd__mux4_2 _14212_ (.A0(\w[57][14] ),
    .A1(\w[61][14] ),
    .A2(\w[59][14] ),
    .A3(\w[63][14] ),
    .S0(net465),
    .S1(net468),
    .X(_03886_));
 sky130_fd_sc_hd__mux4_2 _14213_ (.A0(_03883_),
    .A1(_03884_),
    .A2(_03885_),
    .A3(_03886_),
    .S0(\count16_2[3] ),
    .S1(net454),
    .X(_03887_));
 sky130_fd_sc_hd__mux2i_4 _14214_ (.A0(_03882_),
    .A1(_03887_),
    .S(net453),
    .Y(_11944_));
 sky130_fd_sc_hd__mux4_2 _14215_ (.A0(\w[1][2] ),
    .A1(\w[5][2] ),
    .A2(\w[3][2] ),
    .A3(\w[7][2] ),
    .S0(net422),
    .S1(net429),
    .X(_03888_));
 sky130_fd_sc_hd__mux4_2 _14216_ (.A0(\w[9][2] ),
    .A1(\w[13][2] ),
    .A2(\w[11][2] ),
    .A3(\w[15][2] ),
    .S0(net422),
    .S1(net429),
    .X(_03889_));
 sky130_fd_sc_hd__mux4_2 _14217_ (.A0(\w[17][2] ),
    .A1(\w[21][2] ),
    .A2(\w[19][2] ),
    .A3(\w[23][2] ),
    .S0(net422),
    .S1(net429),
    .X(_03890_));
 sky130_fd_sc_hd__mux4_2 _14218_ (.A0(\w[25][2] ),
    .A1(\w[29][2] ),
    .A2(\w[27][2] ),
    .A3(\w[31][2] ),
    .S0(net422),
    .S1(net429),
    .X(_03891_));
 sky130_fd_sc_hd__mux4_2 _14219_ (.A0(_03888_),
    .A1(_03889_),
    .A2(_03890_),
    .A3(_03891_),
    .S0(net416),
    .S1(net414),
    .X(_03892_));
 sky130_fd_sc_hd__mux4_2 _14220_ (.A0(\w[33][2] ),
    .A1(\w[37][2] ),
    .A2(\w[35][2] ),
    .A3(\w[39][2] ),
    .S0(net423),
    .S1(net427),
    .X(_03893_));
 sky130_fd_sc_hd__mux4_2 _14221_ (.A0(\w[41][2] ),
    .A1(\w[45][2] ),
    .A2(\w[43][2] ),
    .A3(\w[47][2] ),
    .S0(net423),
    .S1(net427),
    .X(_03894_));
 sky130_fd_sc_hd__mux4_2 _14222_ (.A0(\w[49][2] ),
    .A1(\w[53][2] ),
    .A2(\w[51][2] ),
    .A3(\w[55][2] ),
    .S0(net423),
    .S1(net427),
    .X(_03895_));
 sky130_fd_sc_hd__mux4_2 _14223_ (.A0(\w[57][2] ),
    .A1(\w[61][2] ),
    .A2(\w[59][2] ),
    .A3(\w[63][2] ),
    .S0(net423),
    .S1(net427),
    .X(_03896_));
 sky130_fd_sc_hd__mux4_2 _14224_ (.A0(_03893_),
    .A1(_03894_),
    .A2(_03895_),
    .A3(_03896_),
    .S0(net416),
    .S1(net414),
    .X(_03897_));
 sky130_fd_sc_hd__mux2i_4 _14225_ (.A0(_03892_),
    .A1(_03897_),
    .S(net413),
    .Y(_03898_));
 sky130_fd_sc_hd__xnor2_1 _14226_ (.A(_03803_),
    .B(_03898_),
    .Y(_03899_));
 sky130_fd_sc_hd__xnor2_1 _14227_ (.A(_03389_),
    .B(_03899_),
    .Y(_11949_));
 sky130_fd_sc_hd__mux4_2 _14228_ (.A0(\w[0][1] ),
    .A1(\w[4][1] ),
    .A2(\w[2][1] ),
    .A3(\w[6][1] ),
    .S0(net500),
    .S1(net507),
    .X(_03900_));
 sky130_fd_sc_hd__mux4_2 _14229_ (.A0(\w[8][1] ),
    .A1(\w[12][1] ),
    .A2(\w[10][1] ),
    .A3(\w[14][1] ),
    .S0(net500),
    .S1(net507),
    .X(_03901_));
 sky130_fd_sc_hd__mux4_2 _14230_ (.A0(\w[16][1] ),
    .A1(\w[20][1] ),
    .A2(\w[18][1] ),
    .A3(\w[22][1] ),
    .S0(net500),
    .S1(net507),
    .X(_03902_));
 sky130_fd_sc_hd__mux4_2 _14231_ (.A0(\w[24][1] ),
    .A1(\w[28][1] ),
    .A2(\w[26][1] ),
    .A3(\w[30][1] ),
    .S0(net500),
    .S1(net507),
    .X(_03903_));
 sky130_fd_sc_hd__mux4_2 _14232_ (.A0(_03900_),
    .A1(_03901_),
    .A2(_03902_),
    .A3(_03903_),
    .S0(net497),
    .S1(net495),
    .X(_03904_));
 sky130_fd_sc_hd__mux4_2 _14233_ (.A0(\w[32][1] ),
    .A1(\w[36][1] ),
    .A2(\w[34][1] ),
    .A3(\w[38][1] ),
    .S0(net504),
    .S1(net510),
    .X(_03905_));
 sky130_fd_sc_hd__mux4_2 _14234_ (.A0(\w[40][1] ),
    .A1(\w[44][1] ),
    .A2(\w[42][1] ),
    .A3(\w[46][1] ),
    .S0(net504),
    .S1(net510),
    .X(_03906_));
 sky130_fd_sc_hd__mux4_2 _14235_ (.A0(\w[48][1] ),
    .A1(\w[52][1] ),
    .A2(\w[50][1] ),
    .A3(\w[54][1] ),
    .S0(net504),
    .S1(net510),
    .X(_03907_));
 sky130_fd_sc_hd__mux4_2 _14236_ (.A0(\w[56][1] ),
    .A1(\w[60][1] ),
    .A2(\w[58][1] ),
    .A3(\w[62][1] ),
    .S0(net504),
    .S1(net510),
    .X(_03908_));
 sky130_fd_sc_hd__mux4_2 _14237_ (.A0(_03905_),
    .A1(_03906_),
    .A2(_03907_),
    .A3(_03908_),
    .S0(net497),
    .S1(net495),
    .X(_03909_));
 sky130_fd_sc_hd__mux2i_4 _14238_ (.A0(_03904_),
    .A1(_03909_),
    .S(net492),
    .Y(_03910_));
 sky130_fd_sc_hd__xnor2_1 _14239_ (.A(_03264_),
    .B(_03910_),
    .Y(_03911_));
 sky130_fd_sc_hd__xnor2_1 _14240_ (.A(_02853_),
    .B(_03911_),
    .Y(_11948_));
 sky130_fd_sc_hd__mux4_2 _14241_ (.A0(\w[0][15] ),
    .A1(\w[4][15] ),
    .A2(\w[2][15] ),
    .A3(\w[6][15] ),
    .S0(net387),
    .S1(net388),
    .X(_03912_));
 sky130_fd_sc_hd__mux4_2 _14242_ (.A0(\w[8][15] ),
    .A1(\w[12][15] ),
    .A2(\w[10][15] ),
    .A3(\w[14][15] ),
    .S0(net387),
    .S1(net388),
    .X(_03913_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1464 ();
 sky130_fd_sc_hd__mux4_2 _14244_ (.A0(\w[16][15] ),
    .A1(\w[20][15] ),
    .A2(\w[18][15] ),
    .A3(\w[22][15] ),
    .S0(net387),
    .S1(net388),
    .X(_03915_));
 sky130_fd_sc_hd__mux4_2 _14245_ (.A0(\w[24][15] ),
    .A1(\w[28][15] ),
    .A2(\w[26][15] ),
    .A3(\w[30][15] ),
    .S0(net387),
    .S1(net388),
    .X(_03916_));
 sky130_fd_sc_hd__mux4_2 _14246_ (.A0(_03912_),
    .A1(_03913_),
    .A2(_03915_),
    .A3(_03916_),
    .S0(\count7_2[3] ),
    .S1(net376),
    .X(_03917_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1463 ();
 sky130_fd_sc_hd__mux4_2 _14248_ (.A0(\w[32][15] ),
    .A1(\w[36][15] ),
    .A2(\w[34][15] ),
    .A3(\w[38][15] ),
    .S0(net387),
    .S1(\count7_2[1] ),
    .X(_03919_));
 sky130_fd_sc_hd__mux4_2 _14249_ (.A0(\w[40][15] ),
    .A1(\w[44][15] ),
    .A2(\w[42][15] ),
    .A3(\w[46][15] ),
    .S0(net387),
    .S1(net388),
    .X(_03920_));
 sky130_fd_sc_hd__mux4_2 _14250_ (.A0(\w[48][15] ),
    .A1(\w[52][15] ),
    .A2(\w[50][15] ),
    .A3(\w[54][15] ),
    .S0(net387),
    .S1(net388),
    .X(_03921_));
 sky130_fd_sc_hd__mux4_2 _14251_ (.A0(\w[56][15] ),
    .A1(\w[60][15] ),
    .A2(\w[58][15] ),
    .A3(\w[62][15] ),
    .S0(net387),
    .S1(net388),
    .X(_03922_));
 sky130_fd_sc_hd__mux4_2 _14252_ (.A0(_03919_),
    .A1(_03920_),
    .A2(_03921_),
    .A3(_03922_),
    .S0(net379),
    .S1(net376),
    .X(_03923_));
 sky130_fd_sc_hd__mux2i_4 _14253_ (.A0(_03917_),
    .A1(_03923_),
    .S(net373),
    .Y(_11947_));
 sky130_fd_sc_hd__mux4_2 _14254_ (.A0(\w[1][15] ),
    .A1(\w[5][15] ),
    .A2(\w[3][15] ),
    .A3(\w[7][15] ),
    .S0(net466),
    .S1(\count16_2[1] ),
    .X(_03924_));
 sky130_fd_sc_hd__mux4_2 _14255_ (.A0(\w[9][15] ),
    .A1(\w[13][15] ),
    .A2(\w[11][15] ),
    .A3(\w[15][15] ),
    .S0(net466),
    .S1(\count16_2[1] ),
    .X(_03925_));
 sky130_fd_sc_hd__mux4_2 _14256_ (.A0(\w[17][15] ),
    .A1(\w[21][15] ),
    .A2(\w[19][15] ),
    .A3(\w[23][15] ),
    .S0(net466),
    .S1(\count16_2[1] ),
    .X(_03926_));
 sky130_fd_sc_hd__mux4_2 _14257_ (.A0(\w[25][15] ),
    .A1(\w[29][15] ),
    .A2(\w[27][15] ),
    .A3(\w[31][15] ),
    .S0(net466),
    .S1(\count16_2[1] ),
    .X(_03927_));
 sky130_fd_sc_hd__mux4_2 _14258_ (.A0(_03924_),
    .A1(_03925_),
    .A2(_03926_),
    .A3(_03927_),
    .S0(net457),
    .S1(\count16_2[4] ),
    .X(_03928_));
 sky130_fd_sc_hd__mux4_2 _14259_ (.A0(\w[33][15] ),
    .A1(\w[37][15] ),
    .A2(\w[35][15] ),
    .A3(\w[39][15] ),
    .S0(net466),
    .S1(net471),
    .X(_03929_));
 sky130_fd_sc_hd__mux4_2 _14260_ (.A0(\w[41][15] ),
    .A1(\w[45][15] ),
    .A2(\w[43][15] ),
    .A3(\w[47][15] ),
    .S0(net466),
    .S1(net471),
    .X(_03930_));
 sky130_fd_sc_hd__mux4_2 _14261_ (.A0(\w[49][15] ),
    .A1(\w[53][15] ),
    .A2(\w[51][15] ),
    .A3(\w[55][15] ),
    .S0(net466),
    .S1(net471),
    .X(_03931_));
 sky130_fd_sc_hd__mux4_2 _14262_ (.A0(\w[57][15] ),
    .A1(\w[61][15] ),
    .A2(\w[59][15] ),
    .A3(\w[63][15] ),
    .S0(net466),
    .S1(net471),
    .X(_03932_));
 sky130_fd_sc_hd__mux4_2 _14263_ (.A0(_03929_),
    .A1(_03930_),
    .A2(_03931_),
    .A3(_03932_),
    .S0(net457),
    .S1(\count16_2[4] ),
    .X(_03933_));
 sky130_fd_sc_hd__mux2i_4 _14264_ (.A0(_03928_),
    .A1(_03933_),
    .S(\count16_2[5] ),
    .Y(_11952_));
 sky130_fd_sc_hd__mux4_2 _14265_ (.A0(\w[1][3] ),
    .A1(\w[5][3] ),
    .A2(\w[3][3] ),
    .A3(\w[7][3] ),
    .S0(net424),
    .S1(net431),
    .X(_03934_));
 sky130_fd_sc_hd__mux4_2 _14266_ (.A0(\w[9][3] ),
    .A1(\w[13][3] ),
    .A2(\w[11][3] ),
    .A3(\w[15][3] ),
    .S0(net424),
    .S1(net431),
    .X(_03935_));
 sky130_fd_sc_hd__mux4_2 _14267_ (.A0(\w[17][3] ),
    .A1(\w[21][3] ),
    .A2(\w[19][3] ),
    .A3(\w[23][3] ),
    .S0(net424),
    .S1(net431),
    .X(_03936_));
 sky130_fd_sc_hd__mux4_2 _14268_ (.A0(\w[25][3] ),
    .A1(\w[29][3] ),
    .A2(\w[27][3] ),
    .A3(\w[31][3] ),
    .S0(net424),
    .S1(net431),
    .X(_03937_));
 sky130_fd_sc_hd__mux4_2 _14269_ (.A0(_03934_),
    .A1(_03935_),
    .A2(_03936_),
    .A3(_03937_),
    .S0(net417),
    .S1(net540),
    .X(_03938_));
 sky130_fd_sc_hd__mux4_2 _14270_ (.A0(\w[33][3] ),
    .A1(\w[37][3] ),
    .A2(\w[35][3] ),
    .A3(\w[39][3] ),
    .S0(net424),
    .S1(net431),
    .X(_03939_));
 sky130_fd_sc_hd__mux4_2 _14271_ (.A0(\w[41][3] ),
    .A1(\w[45][3] ),
    .A2(\w[43][3] ),
    .A3(\w[47][3] ),
    .S0(net424),
    .S1(net431),
    .X(_03940_));
 sky130_fd_sc_hd__mux4_2 _14272_ (.A0(\w[49][3] ),
    .A1(\w[53][3] ),
    .A2(\w[51][3] ),
    .A3(\w[55][3] ),
    .S0(net424),
    .S1(net431),
    .X(_03941_));
 sky130_fd_sc_hd__mux4_2 _14273_ (.A0(\w[57][3] ),
    .A1(\w[61][3] ),
    .A2(\w[59][3] ),
    .A3(\w[63][3] ),
    .S0(net424),
    .S1(net431),
    .X(_03942_));
 sky130_fd_sc_hd__mux4_2 _14274_ (.A0(_03939_),
    .A1(_03940_),
    .A2(_03941_),
    .A3(_03942_),
    .S0(net417),
    .S1(net540),
    .X(_03943_));
 sky130_fd_sc_hd__mux2i_4 _14275_ (.A0(_03938_),
    .A1(_03943_),
    .S(net413),
    .Y(_03944_));
 sky130_fd_sc_hd__xnor2_1 _14276_ (.A(_03849_),
    .B(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__xnor2_1 _14277_ (.A(_03448_),
    .B(_03945_),
    .Y(_11957_));
 sky130_fd_sc_hd__mux4_2 _14278_ (.A0(\w[0][2] ),
    .A1(\w[4][2] ),
    .A2(\w[2][2] ),
    .A3(\w[6][2] ),
    .S0(net498),
    .S1(net506),
    .X(_03946_));
 sky130_fd_sc_hd__mux4_2 _14279_ (.A0(\w[8][2] ),
    .A1(\w[12][2] ),
    .A2(\w[10][2] ),
    .A3(\w[14][2] ),
    .S0(net498),
    .S1(net506),
    .X(_03947_));
 sky130_fd_sc_hd__mux4_2 _14280_ (.A0(\w[16][2] ),
    .A1(\w[20][2] ),
    .A2(\w[18][2] ),
    .A3(\w[22][2] ),
    .S0(net498),
    .S1(net506),
    .X(_03948_));
 sky130_fd_sc_hd__mux4_2 _14281_ (.A0(\w[24][2] ),
    .A1(\w[28][2] ),
    .A2(\w[26][2] ),
    .A3(\w[30][2] ),
    .S0(net498),
    .S1(net506),
    .X(_03949_));
 sky130_fd_sc_hd__mux4_2 _14282_ (.A0(_03946_),
    .A1(_03947_),
    .A2(_03948_),
    .A3(_03949_),
    .S0(net496),
    .S1(net547),
    .X(_03950_));
 sky130_fd_sc_hd__mux4_2 _14283_ (.A0(\w[32][2] ),
    .A1(\w[36][2] ),
    .A2(\w[34][2] ),
    .A3(\w[38][2] ),
    .S0(net505),
    .S1(net511),
    .X(_03951_));
 sky130_fd_sc_hd__mux4_2 _14284_ (.A0(\w[40][2] ),
    .A1(\w[44][2] ),
    .A2(\w[42][2] ),
    .A3(\w[46][2] ),
    .S0(net505),
    .S1(net511),
    .X(_03952_));
 sky130_fd_sc_hd__mux4_2 _14285_ (.A0(\w[48][2] ),
    .A1(\w[52][2] ),
    .A2(\w[50][2] ),
    .A3(\w[54][2] ),
    .S0(net505),
    .S1(net511),
    .X(_03953_));
 sky130_fd_sc_hd__mux4_2 _14286_ (.A0(\w[56][2] ),
    .A1(\w[60][2] ),
    .A2(\w[58][2] ),
    .A3(\w[62][2] ),
    .S0(net505),
    .S1(net511),
    .X(_03954_));
 sky130_fd_sc_hd__mux4_2 _14287_ (.A0(_03951_),
    .A1(_03952_),
    .A2(_03953_),
    .A3(_03954_),
    .S0(\count15_2[3] ),
    .S1(net547),
    .X(_03955_));
 sky130_fd_sc_hd__mux2i_4 _14288_ (.A0(_03950_),
    .A1(_03955_),
    .S(net493),
    .Y(_03956_));
 sky130_fd_sc_hd__xnor2_1 _14289_ (.A(_03333_),
    .B(_03956_),
    .Y(_03957_));
 sky130_fd_sc_hd__xnor2_1 _14290_ (.A(_03005_),
    .B(_03957_),
    .Y(_11956_));
 sky130_fd_sc_hd__mux4_2 _14291_ (.A0(\w[0][16] ),
    .A1(\w[4][16] ),
    .A2(\w[2][16] ),
    .A3(\w[6][16] ),
    .S0(net387),
    .S1(net388),
    .X(_03958_));
 sky130_fd_sc_hd__mux4_2 _14292_ (.A0(\w[8][16] ),
    .A1(\w[12][16] ),
    .A2(\w[10][16] ),
    .A3(\w[14][16] ),
    .S0(net387),
    .S1(\count7_2[1] ),
    .X(_03959_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1462 ();
 sky130_fd_sc_hd__mux4_2 _14294_ (.A0(\w[16][16] ),
    .A1(\w[20][16] ),
    .A2(\w[18][16] ),
    .A3(\w[22][16] ),
    .S0(net387),
    .S1(\count7_2[1] ),
    .X(_03961_));
 sky130_fd_sc_hd__mux4_2 _14295_ (.A0(\w[24][16] ),
    .A1(\w[28][16] ),
    .A2(\w[26][16] ),
    .A3(\w[30][16] ),
    .S0(net387),
    .S1(net388),
    .X(_03962_));
 sky130_fd_sc_hd__mux4_2 _14296_ (.A0(_03958_),
    .A1(_03959_),
    .A2(_03961_),
    .A3(_03962_),
    .S0(\count7_2[3] ),
    .S1(net376),
    .X(_03963_));
 sky130_fd_sc_hd__mux4_2 _14297_ (.A0(\w[32][16] ),
    .A1(\w[36][16] ),
    .A2(\w[34][16] ),
    .A3(\w[38][16] ),
    .S0(\count7_2[2] ),
    .S1(net393),
    .X(_03964_));
 sky130_fd_sc_hd__mux4_2 _14298_ (.A0(\w[40][16] ),
    .A1(\w[44][16] ),
    .A2(\w[42][16] ),
    .A3(\w[46][16] ),
    .S0(\count7_2[2] ),
    .S1(net393),
    .X(_03965_));
 sky130_fd_sc_hd__mux4_2 _14299_ (.A0(\w[48][16] ),
    .A1(\w[52][16] ),
    .A2(\w[50][16] ),
    .A3(\w[54][16] ),
    .S0(\count7_2[2] ),
    .S1(net393),
    .X(_03966_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1461 ();
 sky130_fd_sc_hd__mux4_2 _14301_ (.A0(\w[56][16] ),
    .A1(\w[60][16] ),
    .A2(\w[58][16] ),
    .A3(\w[62][16] ),
    .S0(\count7_2[2] ),
    .S1(net393),
    .X(_03968_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1460 ();
 sky130_fd_sc_hd__mux4_2 _14303_ (.A0(_03964_),
    .A1(_03965_),
    .A2(_03966_),
    .A3(_03968_),
    .S0(net378),
    .S1(net376),
    .X(_03970_));
 sky130_fd_sc_hd__mux2i_4 _14304_ (.A0(_03963_),
    .A1(_03970_),
    .S(net374),
    .Y(_11955_));
 sky130_fd_sc_hd__mux4_2 _14305_ (.A0(\w[1][16] ),
    .A1(\w[5][16] ),
    .A2(\w[3][16] ),
    .A3(\w[7][16] ),
    .S0(net464),
    .S1(net468),
    .X(_03971_));
 sky130_fd_sc_hd__mux4_2 _14306_ (.A0(\w[9][16] ),
    .A1(\w[13][16] ),
    .A2(\w[11][16] ),
    .A3(\w[15][16] ),
    .S0(net464),
    .S1(net468),
    .X(_03972_));
 sky130_fd_sc_hd__mux4_2 _14307_ (.A0(\w[17][16] ),
    .A1(\w[21][16] ),
    .A2(\w[19][16] ),
    .A3(\w[23][16] ),
    .S0(net464),
    .S1(net468),
    .X(_03973_));
 sky130_fd_sc_hd__mux4_2 _14308_ (.A0(\w[25][16] ),
    .A1(\w[29][16] ),
    .A2(\w[27][16] ),
    .A3(\w[31][16] ),
    .S0(net464),
    .S1(net468),
    .X(_03974_));
 sky130_fd_sc_hd__mux4_2 _14309_ (.A0(_03971_),
    .A1(_03972_),
    .A2(_03973_),
    .A3(_03974_),
    .S0(\count16_2[3] ),
    .S1(net454),
    .X(_03975_));
 sky130_fd_sc_hd__mux4_2 _14310_ (.A0(\w[33][16] ),
    .A1(\w[37][16] ),
    .A2(\w[35][16] ),
    .A3(\w[39][16] ),
    .S0(net465),
    .S1(net469),
    .X(_03976_));
 sky130_fd_sc_hd__mux4_2 _14311_ (.A0(\w[41][16] ),
    .A1(\w[45][16] ),
    .A2(\w[43][16] ),
    .A3(\w[47][16] ),
    .S0(net465),
    .S1(net467),
    .X(_03977_));
 sky130_fd_sc_hd__mux4_2 _14312_ (.A0(\w[49][16] ),
    .A1(\w[53][16] ),
    .A2(\w[51][16] ),
    .A3(\w[55][16] ),
    .S0(net465),
    .S1(net469),
    .X(_03978_));
 sky130_fd_sc_hd__mux4_2 _14313_ (.A0(\w[57][16] ),
    .A1(\w[61][16] ),
    .A2(\w[59][16] ),
    .A3(\w[63][16] ),
    .S0(net465),
    .S1(net469),
    .X(_03979_));
 sky130_fd_sc_hd__mux4_2 _14314_ (.A0(_03976_),
    .A1(_03977_),
    .A2(_03978_),
    .A3(_03979_),
    .S0(\count16_2[3] ),
    .S1(net543),
    .X(_03980_));
 sky130_fd_sc_hd__mux2i_2 _14315_ (.A0(_03975_),
    .A1(_03980_),
    .S(net453),
    .Y(_11960_));
 sky130_fd_sc_hd__mux4_2 _14316_ (.A0(\w[1][4] ),
    .A1(\w[5][4] ),
    .A2(\w[3][4] ),
    .A3(\w[7][4] ),
    .S0(net422),
    .S1(net429),
    .X(_03981_));
 sky130_fd_sc_hd__mux4_2 _14317_ (.A0(\w[9][4] ),
    .A1(\w[13][4] ),
    .A2(\w[11][4] ),
    .A3(\w[15][4] ),
    .S0(net422),
    .S1(net429),
    .X(_03982_));
 sky130_fd_sc_hd__mux4_2 _14318_ (.A0(\w[17][4] ),
    .A1(\w[21][4] ),
    .A2(\w[19][4] ),
    .A3(\w[23][4] ),
    .S0(net422),
    .S1(net429),
    .X(_03983_));
 sky130_fd_sc_hd__mux4_2 _14319_ (.A0(\w[25][4] ),
    .A1(\w[29][4] ),
    .A2(\w[27][4] ),
    .A3(\w[31][4] ),
    .S0(net422),
    .S1(net429),
    .X(_03984_));
 sky130_fd_sc_hd__mux4_2 _14320_ (.A0(_03981_),
    .A1(_03982_),
    .A2(_03983_),
    .A3(_03984_),
    .S0(net416),
    .S1(net414),
    .X(_03985_));
 sky130_fd_sc_hd__mux4_2 _14321_ (.A0(\w[33][4] ),
    .A1(\w[37][4] ),
    .A2(\w[35][4] ),
    .A3(\w[39][4] ),
    .S0(net423),
    .S1(net427),
    .X(_03986_));
 sky130_fd_sc_hd__mux4_2 _14322_ (.A0(\w[41][4] ),
    .A1(\w[45][4] ),
    .A2(\w[43][4] ),
    .A3(\w[47][4] ),
    .S0(net423),
    .S1(net428),
    .X(_03987_));
 sky130_fd_sc_hd__mux4_2 _14323_ (.A0(\w[49][4] ),
    .A1(\w[53][4] ),
    .A2(\w[51][4] ),
    .A3(\w[55][4] ),
    .S0(net423),
    .S1(net428),
    .X(_03988_));
 sky130_fd_sc_hd__mux4_2 _14324_ (.A0(\w[57][4] ),
    .A1(\w[61][4] ),
    .A2(\w[59][4] ),
    .A3(\w[63][4] ),
    .S0(net423),
    .S1(net428),
    .X(_03989_));
 sky130_fd_sc_hd__mux4_2 _14325_ (.A0(_03986_),
    .A1(_03987_),
    .A2(_03988_),
    .A3(_03989_),
    .S0(net417),
    .S1(net414),
    .X(_03990_));
 sky130_fd_sc_hd__mux2i_4 _14326_ (.A0(_03985_),
    .A1(_03990_),
    .S(net413),
    .Y(_03991_));
 sky130_fd_sc_hd__xnor2_1 _14327_ (.A(_03898_),
    .B(_03991_),
    .Y(_03992_));
 sky130_fd_sc_hd__xnor2_1 _14328_ (.A(_03507_),
    .B(_03992_),
    .Y(_11965_));
 sky130_fd_sc_hd__xnor2_1 _14329_ (.A(_03109_),
    .B(_03413_),
    .Y(_03993_));
 sky130_fd_sc_hd__xnor2_1 _14330_ (.A(_02824_),
    .B(_03993_),
    .Y(_11964_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1459 ();
 sky130_fd_sc_hd__mux4_2 _14332_ (.A0(\w[0][17] ),
    .A1(\w[4][17] ),
    .A2(\w[2][17] ),
    .A3(\w[6][17] ),
    .S0(net384),
    .S1(net391),
    .X(_03995_));
 sky130_fd_sc_hd__mux4_2 _14333_ (.A0(\w[8][17] ),
    .A1(\w[12][17] ),
    .A2(\w[10][17] ),
    .A3(\w[14][17] ),
    .S0(net386),
    .S1(net393),
    .X(_03996_));
 sky130_fd_sc_hd__mux4_2 _14334_ (.A0(\w[16][17] ),
    .A1(\w[20][17] ),
    .A2(\w[18][17] ),
    .A3(\w[22][17] ),
    .S0(net384),
    .S1(net391),
    .X(_03997_));
 sky130_fd_sc_hd__mux4_2 _14335_ (.A0(\w[24][17] ),
    .A1(\w[28][17] ),
    .A2(\w[26][17] ),
    .A3(\w[30][17] ),
    .S0(net384),
    .S1(net391),
    .X(_03998_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1458 ();
 sky130_fd_sc_hd__mux4_2 _14337_ (.A0(_03995_),
    .A1(_03996_),
    .A2(_03997_),
    .A3(_03998_),
    .S0(net377),
    .S1(net375),
    .X(_04000_));
 sky130_fd_sc_hd__mux4_2 _14338_ (.A0(\w[32][17] ),
    .A1(\w[36][17] ),
    .A2(\w[34][17] ),
    .A3(\w[38][17] ),
    .S0(net384),
    .S1(net391),
    .X(_04001_));
 sky130_fd_sc_hd__mux4_2 _14339_ (.A0(\w[40][17] ),
    .A1(\w[44][17] ),
    .A2(\w[42][17] ),
    .A3(\w[46][17] ),
    .S0(net384),
    .S1(net391),
    .X(_04002_));
 sky130_fd_sc_hd__mux4_2 _14340_ (.A0(\w[48][17] ),
    .A1(\w[52][17] ),
    .A2(\w[50][17] ),
    .A3(\w[54][17] ),
    .S0(net384),
    .S1(net391),
    .X(_04003_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1457 ();
 sky130_fd_sc_hd__mux4_2 _14342_ (.A0(\w[56][17] ),
    .A1(\w[60][17] ),
    .A2(\w[58][17] ),
    .A3(\w[62][17] ),
    .S0(net384),
    .S1(net391),
    .X(_04005_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1456 ();
 sky130_fd_sc_hd__mux4_2 _14344_ (.A0(_04001_),
    .A1(_04002_),
    .A2(_04003_),
    .A3(_04005_),
    .S0(net377),
    .S1(net375),
    .X(_04007_));
 sky130_fd_sc_hd__mux2i_4 _14345_ (.A0(_04000_),
    .A1(_04007_),
    .S(net373),
    .Y(_11963_));
 sky130_fd_sc_hd__mux4_2 _14346_ (.A0(\w[1][17] ),
    .A1(\w[5][17] ),
    .A2(\w[3][17] ),
    .A3(\w[7][17] ),
    .S0(net459),
    .S1(net470),
    .X(_04008_));
 sky130_fd_sc_hd__mux4_2 _14347_ (.A0(\w[9][17] ),
    .A1(\w[13][17] ),
    .A2(\w[11][17] ),
    .A3(\w[15][17] ),
    .S0(net459),
    .S1(net470),
    .X(_04009_));
 sky130_fd_sc_hd__mux4_2 _14348_ (.A0(\w[17][17] ),
    .A1(\w[21][17] ),
    .A2(\w[19][17] ),
    .A3(\w[23][17] ),
    .S0(net459),
    .S1(net470),
    .X(_04010_));
 sky130_fd_sc_hd__mux4_2 _14349_ (.A0(\w[25][17] ),
    .A1(\w[29][17] ),
    .A2(\w[27][17] ),
    .A3(\w[31][17] ),
    .S0(net459),
    .S1(net470),
    .X(_04011_));
 sky130_fd_sc_hd__mux4_2 _14350_ (.A0(_04008_),
    .A1(_04009_),
    .A2(_04010_),
    .A3(_04011_),
    .S0(net456),
    .S1(net454),
    .X(_04012_));
 sky130_fd_sc_hd__mux4_2 _14351_ (.A0(\w[33][17] ),
    .A1(\w[37][17] ),
    .A2(\w[35][17] ),
    .A3(\w[39][17] ),
    .S0(net459),
    .S1(net470),
    .X(_04013_));
 sky130_fd_sc_hd__mux4_2 _14352_ (.A0(\w[41][17] ),
    .A1(\w[45][17] ),
    .A2(\w[43][17] ),
    .A3(\w[47][17] ),
    .S0(net459),
    .S1(net470),
    .X(_04014_));
 sky130_fd_sc_hd__mux4_2 _14353_ (.A0(\w[49][17] ),
    .A1(\w[53][17] ),
    .A2(\w[51][17] ),
    .A3(\w[55][17] ),
    .S0(net459),
    .S1(net470),
    .X(_04015_));
 sky130_fd_sc_hd__mux4_2 _14354_ (.A0(\w[57][17] ),
    .A1(\w[61][17] ),
    .A2(\w[59][17] ),
    .A3(\w[63][17] ),
    .S0(net459),
    .S1(net470),
    .X(_04016_));
 sky130_fd_sc_hd__mux4_2 _14355_ (.A0(_04013_),
    .A1(_04014_),
    .A2(_04015_),
    .A3(_04016_),
    .S0(net456),
    .S1(net454),
    .X(_04017_));
 sky130_fd_sc_hd__mux2i_4 _14356_ (.A0(_04012_),
    .A1(_04017_),
    .S(net453),
    .Y(_11968_));
 sky130_fd_sc_hd__mux4_2 _14357_ (.A0(\w[1][5] ),
    .A1(\w[5][5] ),
    .A2(\w[3][5] ),
    .A3(\w[7][5] ),
    .S0(net424),
    .S1(net431),
    .X(_04018_));
 sky130_fd_sc_hd__mux4_2 _14358_ (.A0(\w[9][5] ),
    .A1(\w[13][5] ),
    .A2(\w[11][5] ),
    .A3(\w[15][5] ),
    .S0(net424),
    .S1(net431),
    .X(_04019_));
 sky130_fd_sc_hd__mux4_2 _14359_ (.A0(\w[17][5] ),
    .A1(\w[21][5] ),
    .A2(\w[19][5] ),
    .A3(\w[23][5] ),
    .S0(net424),
    .S1(net431),
    .X(_04020_));
 sky130_fd_sc_hd__mux4_2 _14360_ (.A0(\w[25][5] ),
    .A1(\w[29][5] ),
    .A2(\w[27][5] ),
    .A3(\w[31][5] ),
    .S0(net424),
    .S1(net431),
    .X(_04021_));
 sky130_fd_sc_hd__mux4_2 _14361_ (.A0(_04018_),
    .A1(_04019_),
    .A2(_04020_),
    .A3(_04021_),
    .S0(net417),
    .S1(net414),
    .X(_04022_));
 sky130_fd_sc_hd__mux4_2 _14362_ (.A0(\w[33][5] ),
    .A1(\w[37][5] ),
    .A2(\w[35][5] ),
    .A3(\w[39][5] ),
    .S0(net424),
    .S1(net431),
    .X(_04023_));
 sky130_fd_sc_hd__mux4_2 _14363_ (.A0(\w[41][5] ),
    .A1(\w[45][5] ),
    .A2(\w[43][5] ),
    .A3(\w[47][5] ),
    .S0(net424),
    .S1(net431),
    .X(_04024_));
 sky130_fd_sc_hd__mux4_2 _14364_ (.A0(\w[49][5] ),
    .A1(\w[53][5] ),
    .A2(\w[51][5] ),
    .A3(\w[55][5] ),
    .S0(net424),
    .S1(net431),
    .X(_04025_));
 sky130_fd_sc_hd__mux4_2 _14365_ (.A0(\w[57][5] ),
    .A1(\w[61][5] ),
    .A2(\w[59][5] ),
    .A3(\w[63][5] ),
    .S0(net424),
    .S1(net431),
    .X(_04026_));
 sky130_fd_sc_hd__mux4_2 _14366_ (.A0(_04023_),
    .A1(_04024_),
    .A2(_04025_),
    .A3(_04026_),
    .S0(net417),
    .S1(net540),
    .X(_04027_));
 sky130_fd_sc_hd__mux2i_4 _14367_ (.A0(_04022_),
    .A1(_04027_),
    .S(net413),
    .Y(_04028_));
 sky130_fd_sc_hd__xnor2_1 _14368_ (.A(_03944_),
    .B(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__xnor2_2 _14369_ (.A(_03567_),
    .B(_04029_),
    .Y(_11973_));
 sky130_fd_sc_hd__xnor2_1 _14370_ (.A(_03181_),
    .B(_03471_),
    .Y(_04030_));
 sky130_fd_sc_hd__xnor2_2 _14371_ (.A(_02976_),
    .B(_04030_),
    .Y(_11972_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1455 ();
 sky130_fd_sc_hd__mux4_2 _14373_ (.A0(\w[0][18] ),
    .A1(\w[4][18] ),
    .A2(\w[2][18] ),
    .A3(\w[6][18] ),
    .S0(net385),
    .S1(net392),
    .X(_04032_));
 sky130_fd_sc_hd__mux4_2 _14374_ (.A0(\w[8][18] ),
    .A1(\w[12][18] ),
    .A2(\w[10][18] ),
    .A3(\w[14][18] ),
    .S0(net385),
    .S1(net392),
    .X(_04033_));
 sky130_fd_sc_hd__mux4_2 _14375_ (.A0(\w[16][18] ),
    .A1(\w[20][18] ),
    .A2(\w[18][18] ),
    .A3(\w[22][18] ),
    .S0(net385),
    .S1(net392),
    .X(_04034_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1454 ();
 sky130_fd_sc_hd__mux4_2 _14377_ (.A0(\w[24][18] ),
    .A1(\w[28][18] ),
    .A2(\w[26][18] ),
    .A3(\w[30][18] ),
    .S0(net385),
    .S1(net392),
    .X(_04036_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1453 ();
 sky130_fd_sc_hd__mux4_2 _14379_ (.A0(_04032_),
    .A1(_04033_),
    .A2(_04034_),
    .A3(_04036_),
    .S0(net378),
    .S1(net535),
    .X(_04038_));
 sky130_fd_sc_hd__mux4_2 _14380_ (.A0(\w[32][18] ),
    .A1(\w[36][18] ),
    .A2(\w[34][18] ),
    .A3(\w[38][18] ),
    .S0(net385),
    .S1(net392),
    .X(_04039_));
 sky130_fd_sc_hd__mux4_2 _14381_ (.A0(\w[40][18] ),
    .A1(\w[44][18] ),
    .A2(\w[42][18] ),
    .A3(\w[46][18] ),
    .S0(net385),
    .S1(net392),
    .X(_04040_));
 sky130_fd_sc_hd__mux4_2 _14382_ (.A0(\w[48][18] ),
    .A1(\w[52][18] ),
    .A2(\w[50][18] ),
    .A3(\w[54][18] ),
    .S0(net385),
    .S1(net392),
    .X(_04041_));
 sky130_fd_sc_hd__mux4_2 _14383_ (.A0(\w[56][18] ),
    .A1(\w[60][18] ),
    .A2(\w[58][18] ),
    .A3(\w[62][18] ),
    .S0(net385),
    .S1(net392),
    .X(_04042_));
 sky130_fd_sc_hd__mux4_2 _14384_ (.A0(_04039_),
    .A1(_04040_),
    .A2(_04041_),
    .A3(_04042_),
    .S0(net378),
    .S1(net535),
    .X(_04043_));
 sky130_fd_sc_hd__mux2i_4 _14385_ (.A0(_04038_),
    .A1(_04043_),
    .S(net374),
    .Y(_11971_));
 sky130_fd_sc_hd__mux4_2 _14386_ (.A0(\w[1][18] ),
    .A1(\w[5][18] ),
    .A2(\w[3][18] ),
    .A3(\w[7][18] ),
    .S0(net463),
    .S1(net467),
    .X(_04044_));
 sky130_fd_sc_hd__mux4_2 _14387_ (.A0(\w[9][18] ),
    .A1(\w[13][18] ),
    .A2(\w[11][18] ),
    .A3(\w[15][18] ),
    .S0(net463),
    .S1(net467),
    .X(_04045_));
 sky130_fd_sc_hd__mux4_2 _14388_ (.A0(\w[17][18] ),
    .A1(\w[21][18] ),
    .A2(\w[19][18] ),
    .A3(\w[23][18] ),
    .S0(net463),
    .S1(net467),
    .X(_04046_));
 sky130_fd_sc_hd__mux4_2 _14389_ (.A0(\w[25][18] ),
    .A1(\w[29][18] ),
    .A2(\w[27][18] ),
    .A3(\w[31][18] ),
    .S0(net463),
    .S1(net467),
    .X(_04047_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1452 ();
 sky130_fd_sc_hd__mux4_2 _14391_ (.A0(_04044_),
    .A1(_04045_),
    .A2(_04046_),
    .A3(_04047_),
    .S0(net458),
    .S1(net455),
    .X(_04049_));
 sky130_fd_sc_hd__mux4_2 _14392_ (.A0(\w[33][18] ),
    .A1(\w[37][18] ),
    .A2(\w[35][18] ),
    .A3(\w[39][18] ),
    .S0(net463),
    .S1(net469),
    .X(_04050_));
 sky130_fd_sc_hd__mux4_2 _14393_ (.A0(\w[41][18] ),
    .A1(\w[45][18] ),
    .A2(\w[43][18] ),
    .A3(\w[47][18] ),
    .S0(net465),
    .S1(net469),
    .X(_04051_));
 sky130_fd_sc_hd__mux4_2 _14394_ (.A0(\w[49][18] ),
    .A1(\w[53][18] ),
    .A2(\w[51][18] ),
    .A3(\w[55][18] ),
    .S0(net465),
    .S1(net469),
    .X(_04052_));
 sky130_fd_sc_hd__mux4_2 _14395_ (.A0(\w[57][18] ),
    .A1(\w[61][18] ),
    .A2(\w[59][18] ),
    .A3(\w[63][18] ),
    .S0(net465),
    .S1(net469),
    .X(_04053_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1451 ();
 sky130_fd_sc_hd__mux4_2 _14397_ (.A0(_04050_),
    .A1(_04051_),
    .A2(_04052_),
    .A3(_04053_),
    .S0(net458),
    .S1(net455),
    .X(_04055_));
 sky130_fd_sc_hd__mux2i_4 _14398_ (.A0(_04049_),
    .A1(_04055_),
    .S(net542),
    .Y(_11976_));
 sky130_fd_sc_hd__mux4_2 _14399_ (.A0(\w[1][6] ),
    .A1(\w[5][6] ),
    .A2(\w[3][6] ),
    .A3(\w[7][6] ),
    .S0(net420),
    .S1(net427),
    .X(_04056_));
 sky130_fd_sc_hd__mux4_2 _14400_ (.A0(\w[9][6] ),
    .A1(\w[13][6] ),
    .A2(\w[11][6] ),
    .A3(\w[15][6] ),
    .S0(net420),
    .S1(net427),
    .X(_04057_));
 sky130_fd_sc_hd__mux4_2 _14401_ (.A0(\w[17][6] ),
    .A1(\w[21][6] ),
    .A2(\w[19][6] ),
    .A3(\w[23][6] ),
    .S0(net420),
    .S1(net427),
    .X(_04058_));
 sky130_fd_sc_hd__mux4_2 _14402_ (.A0(\w[25][6] ),
    .A1(\w[29][6] ),
    .A2(\w[27][6] ),
    .A3(\w[31][6] ),
    .S0(net420),
    .S1(net427),
    .X(_04059_));
 sky130_fd_sc_hd__mux4_2 _14403_ (.A0(_04056_),
    .A1(_04057_),
    .A2(_04058_),
    .A3(_04059_),
    .S0(net416),
    .S1(net414),
    .X(_04060_));
 sky130_fd_sc_hd__mux4_2 _14404_ (.A0(\w[33][6] ),
    .A1(\w[37][6] ),
    .A2(\w[35][6] ),
    .A3(\w[39][6] ),
    .S0(net419),
    .S1(net426),
    .X(_04061_));
 sky130_fd_sc_hd__mux4_2 _14405_ (.A0(\w[41][6] ),
    .A1(\w[45][6] ),
    .A2(\w[43][6] ),
    .A3(\w[47][6] ),
    .S0(net419),
    .S1(net426),
    .X(_04062_));
 sky130_fd_sc_hd__mux4_2 _14406_ (.A0(\w[49][6] ),
    .A1(\w[53][6] ),
    .A2(\w[51][6] ),
    .A3(\w[55][6] ),
    .S0(net419),
    .S1(net426),
    .X(_04063_));
 sky130_fd_sc_hd__mux4_2 _14407_ (.A0(\w[57][6] ),
    .A1(\w[61][6] ),
    .A2(\w[59][6] ),
    .A3(\w[63][6] ),
    .S0(net419),
    .S1(net426),
    .X(_04064_));
 sky130_fd_sc_hd__mux4_2 _14408_ (.A0(_04061_),
    .A1(_04062_),
    .A2(_04063_),
    .A3(_04064_),
    .S0(net417),
    .S1(net414),
    .X(_04065_));
 sky130_fd_sc_hd__mux2i_4 _14409_ (.A0(_04060_),
    .A1(_04065_),
    .S(net413),
    .Y(_04066_));
 sky130_fd_sc_hd__xnor2_1 _14410_ (.A(_03991_),
    .B(_04066_),
    .Y(_04067_));
 sky130_fd_sc_hd__xnor2_1 _14411_ (.A(_03633_),
    .B(_04067_),
    .Y(_11981_));
 sky130_fd_sc_hd__xnor2_1 _14412_ (.A(_03264_),
    .B(_03530_),
    .Y(_04068_));
 sky130_fd_sc_hd__xnor2_2 _14413_ (.A(_03098_),
    .B(_04068_),
    .Y(_11980_));
 sky130_fd_sc_hd__mux4_2 _14414_ (.A0(\w[0][19] ),
    .A1(\w[4][19] ),
    .A2(\w[2][19] ),
    .A3(\w[6][19] ),
    .S0(net382),
    .S1(net389),
    .X(_04069_));
 sky130_fd_sc_hd__mux4_2 _14415_ (.A0(\w[8][19] ),
    .A1(\w[12][19] ),
    .A2(\w[10][19] ),
    .A3(\w[14][19] ),
    .S0(net382),
    .S1(net389),
    .X(_04070_));
 sky130_fd_sc_hd__mux4_2 _14416_ (.A0(\w[16][19] ),
    .A1(\w[20][19] ),
    .A2(\w[18][19] ),
    .A3(\w[22][19] ),
    .S0(net382),
    .S1(net389),
    .X(_04071_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1450 ();
 sky130_fd_sc_hd__mux4_2 _14418_ (.A0(\w[24][19] ),
    .A1(\w[28][19] ),
    .A2(\w[26][19] ),
    .A3(\w[30][19] ),
    .S0(net382),
    .S1(net389),
    .X(_04073_));
 sky130_fd_sc_hd__mux4_2 _14419_ (.A0(_04069_),
    .A1(_04070_),
    .A2(_04071_),
    .A3(_04073_),
    .S0(net377),
    .S1(net375),
    .X(_04074_));
 sky130_fd_sc_hd__mux4_2 _14420_ (.A0(\w[32][19] ),
    .A1(\w[36][19] ),
    .A2(\w[34][19] ),
    .A3(\w[38][19] ),
    .S0(net383),
    .S1(net390),
    .X(_04075_));
 sky130_fd_sc_hd__mux4_2 _14421_ (.A0(\w[40][19] ),
    .A1(\w[44][19] ),
    .A2(\w[42][19] ),
    .A3(\w[46][19] ),
    .S0(net383),
    .S1(net390),
    .X(_04076_));
 sky130_fd_sc_hd__mux4_2 _14422_ (.A0(\w[48][19] ),
    .A1(\w[52][19] ),
    .A2(\w[50][19] ),
    .A3(\w[54][19] ),
    .S0(net383),
    .S1(net390),
    .X(_04077_));
 sky130_fd_sc_hd__mux4_2 _14423_ (.A0(\w[56][19] ),
    .A1(\w[60][19] ),
    .A2(\w[58][19] ),
    .A3(\w[62][19] ),
    .S0(net383),
    .S1(net390),
    .X(_04078_));
 sky130_fd_sc_hd__mux4_2 _14424_ (.A0(_04075_),
    .A1(_04076_),
    .A2(_04077_),
    .A3(_04078_),
    .S0(net378),
    .S1(net535),
    .X(_04079_));
 sky130_fd_sc_hd__mux2i_4 _14425_ (.A0(_04074_),
    .A1(_04079_),
    .S(net374),
    .Y(_11979_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1449 ();
 sky130_fd_sc_hd__mux4_2 _14427_ (.A0(\w[1][19] ),
    .A1(\w[5][19] ),
    .A2(\w[3][19] ),
    .A3(\w[7][19] ),
    .S0(net463),
    .S1(net467),
    .X(_04081_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1448 ();
 sky130_fd_sc_hd__mux4_2 _14429_ (.A0(\w[9][19] ),
    .A1(\w[13][19] ),
    .A2(\w[11][19] ),
    .A3(\w[15][19] ),
    .S0(net463),
    .S1(net467),
    .X(_04083_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1447 ();
 sky130_fd_sc_hd__mux4_2 _14431_ (.A0(\w[17][19] ),
    .A1(\w[21][19] ),
    .A2(\w[19][19] ),
    .A3(\w[23][19] ),
    .S0(net463),
    .S1(net467),
    .X(_04085_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1446 ();
 sky130_fd_sc_hd__mux4_2 _14433_ (.A0(\w[25][19] ),
    .A1(\w[29][19] ),
    .A2(\w[27][19] ),
    .A3(\w[31][19] ),
    .S0(net463),
    .S1(net467),
    .X(_04087_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1445 ();
 sky130_fd_sc_hd__mux4_2 _14435_ (.A0(_04081_),
    .A1(_04083_),
    .A2(_04085_),
    .A3(_04087_),
    .S0(net458),
    .S1(net455),
    .X(_04089_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1444 ();
 sky130_fd_sc_hd__mux4_2 _14437_ (.A0(\w[33][19] ),
    .A1(\w[37][19] ),
    .A2(\w[35][19] ),
    .A3(\w[39][19] ),
    .S0(\count16_2[2] ),
    .S1(net469),
    .X(_04091_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1443 ();
 sky130_fd_sc_hd__mux4_2 _14439_ (.A0(\w[41][19] ),
    .A1(\w[45][19] ),
    .A2(\w[43][19] ),
    .A3(\w[47][19] ),
    .S0(\count16_2[2] ),
    .S1(net469),
    .X(_04093_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1442 ();
 sky130_fd_sc_hd__mux4_2 _14441_ (.A0(\w[49][19] ),
    .A1(\w[53][19] ),
    .A2(\w[51][19] ),
    .A3(\w[55][19] ),
    .S0(\count16_2[2] ),
    .S1(net469),
    .X(_04095_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1441 ();
 sky130_fd_sc_hd__mux4_2 _14443_ (.A0(\w[57][19] ),
    .A1(\w[61][19] ),
    .A2(\w[59][19] ),
    .A3(\w[63][19] ),
    .S0(\count16_2[2] ),
    .S1(net469),
    .X(_04097_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1440 ();
 sky130_fd_sc_hd__mux4_2 _14445_ (.A0(_04091_),
    .A1(_04093_),
    .A2(_04095_),
    .A3(_04097_),
    .S0(net458),
    .S1(net455),
    .X(_04099_));
 sky130_fd_sc_hd__mux2i_2 _14446_ (.A0(_04089_),
    .A1(_04099_),
    .S(net542),
    .Y(_11984_));
 sky130_fd_sc_hd__mux4_2 _14447_ (.A0(\w[1][7] ),
    .A1(\w[5][7] ),
    .A2(\w[3][7] ),
    .A3(\w[7][7] ),
    .S0(net424),
    .S1(net431),
    .X(_04100_));
 sky130_fd_sc_hd__mux4_2 _14448_ (.A0(\w[9][7] ),
    .A1(\w[13][7] ),
    .A2(\w[11][7] ),
    .A3(\w[15][7] ),
    .S0(net424),
    .S1(net431),
    .X(_04101_));
 sky130_fd_sc_hd__mux4_2 _14449_ (.A0(\w[17][7] ),
    .A1(\w[21][7] ),
    .A2(\w[19][7] ),
    .A3(\w[23][7] ),
    .S0(net424),
    .S1(net431),
    .X(_04102_));
 sky130_fd_sc_hd__mux4_2 _14450_ (.A0(\w[25][7] ),
    .A1(\w[29][7] ),
    .A2(\w[27][7] ),
    .A3(\w[31][7] ),
    .S0(net424),
    .S1(net431),
    .X(_04103_));
 sky130_fd_sc_hd__mux4_2 _14451_ (.A0(_04100_),
    .A1(_04101_),
    .A2(_04102_),
    .A3(_04103_),
    .S0(\count2_2[3] ),
    .S1(net540),
    .X(_04104_));
 sky130_fd_sc_hd__mux4_2 _14452_ (.A0(\w[33][7] ),
    .A1(\w[37][7] ),
    .A2(\w[35][7] ),
    .A3(\w[39][7] ),
    .S0(net424),
    .S1(net429),
    .X(_04105_));
 sky130_fd_sc_hd__mux4_2 _14453_ (.A0(\w[41][7] ),
    .A1(\w[45][7] ),
    .A2(\w[43][7] ),
    .A3(\w[47][7] ),
    .S0(net424),
    .S1(net429),
    .X(_04106_));
 sky130_fd_sc_hd__mux4_2 _14454_ (.A0(\w[49][7] ),
    .A1(\w[53][7] ),
    .A2(\w[51][7] ),
    .A3(\w[55][7] ),
    .S0(net424),
    .S1(net429),
    .X(_04107_));
 sky130_fd_sc_hd__mux4_2 _14455_ (.A0(\w[57][7] ),
    .A1(\w[61][7] ),
    .A2(\w[59][7] ),
    .A3(\w[63][7] ),
    .S0(net424),
    .S1(net429),
    .X(_04108_));
 sky130_fd_sc_hd__mux4_2 _14456_ (.A0(_04105_),
    .A1(_04106_),
    .A2(_04107_),
    .A3(_04108_),
    .S0(net417),
    .S1(net540),
    .X(_04109_));
 sky130_fd_sc_hd__mux2i_4 _14457_ (.A0(_04104_),
    .A1(_04109_),
    .S(net413),
    .Y(_04110_));
 sky130_fd_sc_hd__xnor2_1 _14458_ (.A(_04028_),
    .B(_04110_),
    .Y(_04111_));
 sky130_fd_sc_hd__xnor2_1 _14459_ (.A(_03697_),
    .B(_04111_),
    .Y(_11989_));
 sky130_fd_sc_hd__xnor2_1 _14460_ (.A(_03333_),
    .B(_03590_),
    .Y(_04112_));
 sky130_fd_sc_hd__xnor2_2 _14461_ (.A(_03194_),
    .B(_04112_),
    .Y(_11988_));
 sky130_fd_sc_hd__mux4_2 _14462_ (.A0(\w[0][20] ),
    .A1(\w[4][20] ),
    .A2(\w[2][20] ),
    .A3(\w[6][20] ),
    .S0(net383),
    .S1(net390),
    .X(_04113_));
 sky130_fd_sc_hd__mux4_2 _14463_ (.A0(\w[8][20] ),
    .A1(\w[12][20] ),
    .A2(\w[10][20] ),
    .A3(\w[14][20] ),
    .S0(net383),
    .S1(net390),
    .X(_04114_));
 sky130_fd_sc_hd__mux4_2 _14464_ (.A0(\w[16][20] ),
    .A1(\w[20][20] ),
    .A2(\w[18][20] ),
    .A3(\w[22][20] ),
    .S0(net383),
    .S1(net390),
    .X(_04115_));
 sky130_fd_sc_hd__mux4_2 _14465_ (.A0(\w[24][20] ),
    .A1(\w[28][20] ),
    .A2(\w[26][20] ),
    .A3(\w[30][20] ),
    .S0(net383),
    .S1(net390),
    .X(_04116_));
 sky130_fd_sc_hd__mux4_2 _14466_ (.A0(_04113_),
    .A1(_04114_),
    .A2(_04115_),
    .A3(_04116_),
    .S0(net378),
    .S1(net535),
    .X(_04117_));
 sky130_fd_sc_hd__mux4_2 _14467_ (.A0(\w[32][20] ),
    .A1(\w[36][20] ),
    .A2(\w[34][20] ),
    .A3(\w[38][20] ),
    .S0(net385),
    .S1(net392),
    .X(_04118_));
 sky130_fd_sc_hd__mux4_2 _14468_ (.A0(\w[40][20] ),
    .A1(\w[44][20] ),
    .A2(\w[42][20] ),
    .A3(\w[46][20] ),
    .S0(net385),
    .S1(net392),
    .X(_04119_));
 sky130_fd_sc_hd__mux4_2 _14469_ (.A0(\w[48][20] ),
    .A1(\w[52][20] ),
    .A2(\w[50][20] ),
    .A3(\w[54][20] ),
    .S0(net385),
    .S1(net392),
    .X(_04120_));
 sky130_fd_sc_hd__mux4_2 _14470_ (.A0(\w[56][20] ),
    .A1(\w[60][20] ),
    .A2(\w[58][20] ),
    .A3(\w[62][20] ),
    .S0(net385),
    .S1(net392),
    .X(_04121_));
 sky130_fd_sc_hd__mux4_2 _14471_ (.A0(_04118_),
    .A1(_04119_),
    .A2(_04120_),
    .A3(_04121_),
    .S0(net378),
    .S1(net535),
    .X(_04122_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1439 ();
 sky130_fd_sc_hd__mux2i_4 _14473_ (.A0(_04117_),
    .A1(_04122_),
    .S(net374),
    .Y(_11987_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1438 ();
 sky130_fd_sc_hd__mux4_2 _14475_ (.A0(\w[1][20] ),
    .A1(\w[5][20] ),
    .A2(\w[3][20] ),
    .A3(\w[7][20] ),
    .S0(net463),
    .S1(net469),
    .X(_04125_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1437 ();
 sky130_fd_sc_hd__mux4_2 _14477_ (.A0(\w[9][20] ),
    .A1(\w[13][20] ),
    .A2(\w[11][20] ),
    .A3(\w[15][20] ),
    .S0(net463),
    .S1(net469),
    .X(_04127_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1436 ();
 sky130_fd_sc_hd__mux4_2 _14479_ (.A0(\w[17][20] ),
    .A1(\w[21][20] ),
    .A2(\w[19][20] ),
    .A3(\w[23][20] ),
    .S0(net463),
    .S1(net469),
    .X(_04129_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1435 ();
 sky130_fd_sc_hd__mux4_2 _14481_ (.A0(\w[25][20] ),
    .A1(\w[29][20] ),
    .A2(\w[27][20] ),
    .A3(\w[31][20] ),
    .S0(net463),
    .S1(net469),
    .X(_04131_));
 sky130_fd_sc_hd__mux4_2 _14482_ (.A0(_04125_),
    .A1(_04127_),
    .A2(_04129_),
    .A3(_04131_),
    .S0(net458),
    .S1(net455),
    .X(_04132_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1434 ();
 sky130_fd_sc_hd__mux4_2 _14484_ (.A0(\w[33][20] ),
    .A1(\w[37][20] ),
    .A2(\w[35][20] ),
    .A3(\w[39][20] ),
    .S0(\count16_2[2] ),
    .S1(net471),
    .X(_04134_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1433 ();
 sky130_fd_sc_hd__mux4_2 _14486_ (.A0(\w[41][20] ),
    .A1(\w[45][20] ),
    .A2(\w[43][20] ),
    .A3(\w[47][20] ),
    .S0(\count16_2[2] ),
    .S1(net471),
    .X(_04136_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1432 ();
 sky130_fd_sc_hd__mux4_2 _14488_ (.A0(\w[49][20] ),
    .A1(\w[53][20] ),
    .A2(\w[51][20] ),
    .A3(\w[55][20] ),
    .S0(\count16_2[2] ),
    .S1(net471),
    .X(_04138_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1431 ();
 sky130_fd_sc_hd__mux4_2 _14490_ (.A0(\w[57][20] ),
    .A1(\w[61][20] ),
    .A2(\w[59][20] ),
    .A3(\w[63][20] ),
    .S0(\count16_2[2] ),
    .S1(net471),
    .X(_04140_));
 sky130_fd_sc_hd__mux4_2 _14491_ (.A0(_04134_),
    .A1(_04136_),
    .A2(_04138_),
    .A3(_04140_),
    .S0(net458),
    .S1(net455),
    .X(_04141_));
 sky130_fd_sc_hd__mux2i_2 _14492_ (.A0(_04132_),
    .A1(_04141_),
    .S(net542),
    .Y(_11992_));
 sky130_fd_sc_hd__mux4_2 _14493_ (.A0(\w[1][8] ),
    .A1(\w[5][8] ),
    .A2(\w[3][8] ),
    .A3(\w[7][8] ),
    .S0(net420),
    .S1(net427),
    .X(_04142_));
 sky130_fd_sc_hd__mux4_2 _14494_ (.A0(\w[9][8] ),
    .A1(\w[13][8] ),
    .A2(\w[11][8] ),
    .A3(\w[15][8] ),
    .S0(net420),
    .S1(net427),
    .X(_04143_));
 sky130_fd_sc_hd__mux4_2 _14495_ (.A0(\w[17][8] ),
    .A1(\w[21][8] ),
    .A2(\w[19][8] ),
    .A3(\w[23][8] ),
    .S0(net420),
    .S1(net427),
    .X(_04144_));
 sky130_fd_sc_hd__mux4_2 _14496_ (.A0(\w[25][8] ),
    .A1(\w[29][8] ),
    .A2(\w[27][8] ),
    .A3(\w[31][8] ),
    .S0(net420),
    .S1(net427),
    .X(_04145_));
 sky130_fd_sc_hd__mux4_2 _14497_ (.A0(_04142_),
    .A1(_04143_),
    .A2(_04144_),
    .A3(_04145_),
    .S0(net416),
    .S1(net414),
    .X(_04146_));
 sky130_fd_sc_hd__mux4_2 _14498_ (.A0(\w[33][8] ),
    .A1(\w[37][8] ),
    .A2(\w[35][8] ),
    .A3(\w[39][8] ),
    .S0(net419),
    .S1(net426),
    .X(_04147_));
 sky130_fd_sc_hd__mux4_2 _14499_ (.A0(\w[41][8] ),
    .A1(\w[45][8] ),
    .A2(\w[43][8] ),
    .A3(\w[47][8] ),
    .S0(net419),
    .S1(net426),
    .X(_04148_));
 sky130_fd_sc_hd__mux4_2 _14500_ (.A0(\w[49][8] ),
    .A1(\w[53][8] ),
    .A2(\w[51][8] ),
    .A3(\w[55][8] ),
    .S0(net419),
    .S1(net426),
    .X(_04149_));
 sky130_fd_sc_hd__mux4_2 _14501_ (.A0(\w[57][8] ),
    .A1(\w[61][8] ),
    .A2(\w[59][8] ),
    .A3(\w[63][8] ),
    .S0(net419),
    .S1(net426),
    .X(_04150_));
 sky130_fd_sc_hd__mux4_2 _14502_ (.A0(_04147_),
    .A1(_04148_),
    .A2(_04149_),
    .A3(_04150_),
    .S0(net417),
    .S1(net415),
    .X(_04151_));
 sky130_fd_sc_hd__mux2i_4 _14503_ (.A0(_04146_),
    .A1(_04151_),
    .S(net413),
    .Y(_04152_));
 sky130_fd_sc_hd__xnor2_1 _14504_ (.A(_04066_),
    .B(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__xnor2_1 _14505_ (.A(_03743_),
    .B(_04153_),
    .Y(_11997_));
 sky130_fd_sc_hd__xnor2_1 _14506_ (.A(_03413_),
    .B(_03645_),
    .Y(_04154_));
 sky130_fd_sc_hd__xnor2_2 _14507_ (.A(_02882_),
    .B(_04154_),
    .Y(_11996_));
 sky130_fd_sc_hd__mux4_2 _14508_ (.A0(\w[0][21] ),
    .A1(\w[4][21] ),
    .A2(\w[2][21] ),
    .A3(\w[6][21] ),
    .S0(net382),
    .S1(net389),
    .X(_04155_));
 sky130_fd_sc_hd__mux4_2 _14509_ (.A0(\w[8][21] ),
    .A1(\w[12][21] ),
    .A2(\w[10][21] ),
    .A3(\w[14][21] ),
    .S0(net382),
    .S1(net389),
    .X(_04156_));
 sky130_fd_sc_hd__mux4_2 _14510_ (.A0(\w[16][21] ),
    .A1(\w[20][21] ),
    .A2(\w[18][21] ),
    .A3(\w[22][21] ),
    .S0(net382),
    .S1(net389),
    .X(_04157_));
 sky130_fd_sc_hd__mux4_2 _14511_ (.A0(\w[24][21] ),
    .A1(\w[28][21] ),
    .A2(\w[26][21] ),
    .A3(\w[30][21] ),
    .S0(net382),
    .S1(net389),
    .X(_04158_));
 sky130_fd_sc_hd__mux4_2 _14512_ (.A0(_04155_),
    .A1(_04156_),
    .A2(_04157_),
    .A3(_04158_),
    .S0(net377),
    .S1(net375),
    .X(_04159_));
 sky130_fd_sc_hd__mux4_2 _14513_ (.A0(\w[32][21] ),
    .A1(\w[36][21] ),
    .A2(\w[34][21] ),
    .A3(\w[38][21] ),
    .S0(net385),
    .S1(net392),
    .X(_04160_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1430 ();
 sky130_fd_sc_hd__mux4_2 _14515_ (.A0(\w[40][21] ),
    .A1(\w[44][21] ),
    .A2(\w[42][21] ),
    .A3(\w[46][21] ),
    .S0(net385),
    .S1(net392),
    .X(_04162_));
 sky130_fd_sc_hd__mux4_2 _14516_ (.A0(\w[48][21] ),
    .A1(\w[52][21] ),
    .A2(\w[50][21] ),
    .A3(\w[54][21] ),
    .S0(net385),
    .S1(net392),
    .X(_04163_));
 sky130_fd_sc_hd__mux4_2 _14517_ (.A0(\w[56][21] ),
    .A1(\w[60][21] ),
    .A2(\w[58][21] ),
    .A3(\w[62][21] ),
    .S0(net385),
    .S1(net392),
    .X(_04164_));
 sky130_fd_sc_hd__mux4_2 _14518_ (.A0(_04160_),
    .A1(_04162_),
    .A2(_04163_),
    .A3(_04164_),
    .S0(net378),
    .S1(\count7_2[4] ),
    .X(_04165_));
 sky130_fd_sc_hd__mux2i_4 _14519_ (.A0(_04159_),
    .A1(_04165_),
    .S(net374),
    .Y(_11995_));
 sky130_fd_sc_hd__mux4_2 _14520_ (.A0(\w[1][21] ),
    .A1(\w[5][21] ),
    .A2(\w[3][21] ),
    .A3(\w[7][21] ),
    .S0(net463),
    .S1(net468),
    .X(_04166_));
 sky130_fd_sc_hd__mux4_2 _14521_ (.A0(\w[9][21] ),
    .A1(\w[13][21] ),
    .A2(\w[11][21] ),
    .A3(\w[15][21] ),
    .S0(net463),
    .S1(net468),
    .X(_04167_));
 sky130_fd_sc_hd__mux4_2 _14522_ (.A0(\w[17][21] ),
    .A1(\w[21][21] ),
    .A2(\w[19][21] ),
    .A3(\w[23][21] ),
    .S0(net463),
    .S1(net467),
    .X(_04168_));
 sky130_fd_sc_hd__mux4_2 _14523_ (.A0(\w[25][21] ),
    .A1(\w[29][21] ),
    .A2(\w[27][21] ),
    .A3(\w[31][21] ),
    .S0(net463),
    .S1(net467),
    .X(_04169_));
 sky130_fd_sc_hd__mux4_2 _14524_ (.A0(_04166_),
    .A1(_04167_),
    .A2(_04168_),
    .A3(_04169_),
    .S0(net458),
    .S1(net455),
    .X(_04170_));
 sky130_fd_sc_hd__mux4_2 _14525_ (.A0(\w[33][21] ),
    .A1(\w[37][21] ),
    .A2(\w[35][21] ),
    .A3(\w[39][21] ),
    .S0(net465),
    .S1(net467),
    .X(_04171_));
 sky130_fd_sc_hd__mux4_2 _14526_ (.A0(\w[41][21] ),
    .A1(\w[45][21] ),
    .A2(\w[43][21] ),
    .A3(\w[47][21] ),
    .S0(net465),
    .S1(net467),
    .X(_04172_));
 sky130_fd_sc_hd__mux4_2 _14527_ (.A0(\w[49][21] ),
    .A1(\w[53][21] ),
    .A2(\w[51][21] ),
    .A3(\w[55][21] ),
    .S0(net465),
    .S1(net467),
    .X(_04173_));
 sky130_fd_sc_hd__mux4_2 _14528_ (.A0(\w[57][21] ),
    .A1(\w[61][21] ),
    .A2(\w[59][21] ),
    .A3(\w[63][21] ),
    .S0(net465),
    .S1(net467),
    .X(_04174_));
 sky130_fd_sc_hd__mux4_2 _14529_ (.A0(_04171_),
    .A1(_04172_),
    .A2(_04173_),
    .A3(_04174_),
    .S0(net458),
    .S1(net455),
    .X(_04175_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1429 ();
 sky130_fd_sc_hd__mux2i_4 _14531_ (.A0(_04170_),
    .A1(_04175_),
    .S(net542),
    .Y(_12000_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1428 ();
 sky130_fd_sc_hd__mux4_2 _14533_ (.A0(\w[1][9] ),
    .A1(\w[5][9] ),
    .A2(\w[3][9] ),
    .A3(\w[7][9] ),
    .S0(net541),
    .S1(net431),
    .X(_04178_));
 sky130_fd_sc_hd__mux4_2 _14534_ (.A0(\w[9][9] ),
    .A1(\w[13][9] ),
    .A2(\w[11][9] ),
    .A3(\w[15][9] ),
    .S0(net541),
    .S1(net431),
    .X(_04179_));
 sky130_fd_sc_hd__mux4_2 _14535_ (.A0(\w[17][9] ),
    .A1(\w[21][9] ),
    .A2(\w[19][9] ),
    .A3(\w[23][9] ),
    .S0(net541),
    .S1(net431),
    .X(_04180_));
 sky130_fd_sc_hd__mux4_2 _14536_ (.A0(\w[25][9] ),
    .A1(\w[29][9] ),
    .A2(\w[27][9] ),
    .A3(\w[31][9] ),
    .S0(net541),
    .S1(net431),
    .X(_04181_));
 sky130_fd_sc_hd__mux4_2 _14537_ (.A0(_04178_),
    .A1(_04179_),
    .A2(_04180_),
    .A3(_04181_),
    .S0(\count2_2[3] ),
    .S1(net540),
    .X(_04182_));
 sky130_fd_sc_hd__mux4_2 _14538_ (.A0(\w[33][9] ),
    .A1(\w[37][9] ),
    .A2(\w[35][9] ),
    .A3(\w[39][9] ),
    .S0(net425),
    .S1(net430),
    .X(_04183_));
 sky130_fd_sc_hd__mux4_2 _14539_ (.A0(\w[41][9] ),
    .A1(\w[45][9] ),
    .A2(\w[43][9] ),
    .A3(\w[47][9] ),
    .S0(net425),
    .S1(net430),
    .X(_04184_));
 sky130_fd_sc_hd__mux4_2 _14540_ (.A0(\w[49][9] ),
    .A1(\w[53][9] ),
    .A2(\w[51][9] ),
    .A3(\w[55][9] ),
    .S0(net425),
    .S1(net430),
    .X(_04185_));
 sky130_fd_sc_hd__mux4_2 _14541_ (.A0(\w[57][9] ),
    .A1(\w[61][9] ),
    .A2(\w[59][9] ),
    .A3(\w[63][9] ),
    .S0(net425),
    .S1(net430),
    .X(_04186_));
 sky130_fd_sc_hd__mux4_2 _14542_ (.A0(_04183_),
    .A1(_04184_),
    .A2(_04185_),
    .A3(_04186_),
    .S0(net417),
    .S1(net414),
    .X(_04187_));
 sky130_fd_sc_hd__mux2i_2 _14543_ (.A0(_04182_),
    .A1(_04187_),
    .S(net539),
    .Y(_04188_));
 sky130_fd_sc_hd__xnor2_1 _14544_ (.A(_04110_),
    .B(_04188_),
    .Y(_12005_));
 sky130_fd_sc_hd__xnor2_1 _14545_ (.A(_03471_),
    .B(_03709_),
    .Y(_04189_));
 sky130_fd_sc_hd__xnor2_1 _14546_ (.A(_02994_),
    .B(_04189_),
    .Y(_12004_));
 sky130_fd_sc_hd__mux4_2 _14547_ (.A0(\w[0][22] ),
    .A1(\w[4][22] ),
    .A2(\w[2][22] ),
    .A3(\w[6][22] ),
    .S0(net381),
    .S1(net389),
    .X(_04190_));
 sky130_fd_sc_hd__mux4_2 _14548_ (.A0(\w[8][22] ),
    .A1(\w[12][22] ),
    .A2(\w[10][22] ),
    .A3(\w[14][22] ),
    .S0(net382),
    .S1(net389),
    .X(_04191_));
 sky130_fd_sc_hd__mux4_2 _14549_ (.A0(\w[16][22] ),
    .A1(\w[20][22] ),
    .A2(\w[18][22] ),
    .A3(\w[22][22] ),
    .S0(net382),
    .S1(net389),
    .X(_04192_));
 sky130_fd_sc_hd__mux4_2 _14550_ (.A0(\w[24][22] ),
    .A1(\w[28][22] ),
    .A2(\w[26][22] ),
    .A3(\w[30][22] ),
    .S0(net382),
    .S1(net389),
    .X(_04193_));
 sky130_fd_sc_hd__mux4_2 _14551_ (.A0(_04190_),
    .A1(_04191_),
    .A2(_04192_),
    .A3(_04193_),
    .S0(net377),
    .S1(net535),
    .X(_04194_));
 sky130_fd_sc_hd__mux4_2 _14552_ (.A0(\w[32][22] ),
    .A1(\w[36][22] ),
    .A2(\w[34][22] ),
    .A3(\w[38][22] ),
    .S0(net381),
    .S1(net389),
    .X(_04195_));
 sky130_fd_sc_hd__mux4_2 _14553_ (.A0(\w[40][22] ),
    .A1(\w[44][22] ),
    .A2(\w[42][22] ),
    .A3(\w[46][22] ),
    .S0(net381),
    .S1(net389),
    .X(_04196_));
 sky130_fd_sc_hd__mux4_2 _14554_ (.A0(\w[48][22] ),
    .A1(\w[52][22] ),
    .A2(\w[50][22] ),
    .A3(\w[54][22] ),
    .S0(net381),
    .S1(net389),
    .X(_04197_));
 sky130_fd_sc_hd__mux4_2 _14555_ (.A0(\w[56][22] ),
    .A1(\w[60][22] ),
    .A2(\w[58][22] ),
    .A3(\w[62][22] ),
    .S0(net381),
    .S1(net389),
    .X(_04198_));
 sky130_fd_sc_hd__mux4_2 _14556_ (.A0(_04195_),
    .A1(_04196_),
    .A2(_04197_),
    .A3(_04198_),
    .S0(net378),
    .S1(net535),
    .X(_04199_));
 sky130_fd_sc_hd__mux2i_4 _14557_ (.A0(_04194_),
    .A1(_04199_),
    .S(net374),
    .Y(_12003_));
 sky130_fd_sc_hd__mux4_2 _14558_ (.A0(\w[1][22] ),
    .A1(\w[5][22] ),
    .A2(\w[3][22] ),
    .A3(\w[7][22] ),
    .S0(net463),
    .S1(net468),
    .X(_04200_));
 sky130_fd_sc_hd__mux4_2 _14559_ (.A0(\w[9][22] ),
    .A1(\w[13][22] ),
    .A2(\w[11][22] ),
    .A3(\w[15][22] ),
    .S0(net463),
    .S1(net468),
    .X(_04201_));
 sky130_fd_sc_hd__mux4_2 _14560_ (.A0(\w[17][22] ),
    .A1(\w[21][22] ),
    .A2(\w[19][22] ),
    .A3(\w[23][22] ),
    .S0(net463),
    .S1(net468),
    .X(_04202_));
 sky130_fd_sc_hd__mux4_2 _14561_ (.A0(\w[25][22] ),
    .A1(\w[29][22] ),
    .A2(\w[27][22] ),
    .A3(\w[31][22] ),
    .S0(net463),
    .S1(net468),
    .X(_04203_));
 sky130_fd_sc_hd__mux4_2 _14562_ (.A0(_04200_),
    .A1(_04201_),
    .A2(_04202_),
    .A3(_04203_),
    .S0(net458),
    .S1(net455),
    .X(_04204_));
 sky130_fd_sc_hd__mux4_2 _14563_ (.A0(\w[33][22] ),
    .A1(\w[37][22] ),
    .A2(\w[35][22] ),
    .A3(\w[39][22] ),
    .S0(net465),
    .S1(net468),
    .X(_04205_));
 sky130_fd_sc_hd__mux4_2 _14564_ (.A0(\w[41][22] ),
    .A1(\w[45][22] ),
    .A2(\w[43][22] ),
    .A3(\w[47][22] ),
    .S0(net465),
    .S1(net468),
    .X(_04206_));
 sky130_fd_sc_hd__mux4_2 _14565_ (.A0(\w[49][22] ),
    .A1(\w[53][22] ),
    .A2(\w[51][22] ),
    .A3(\w[55][22] ),
    .S0(net465),
    .S1(net468),
    .X(_04207_));
 sky130_fd_sc_hd__mux4_2 _14566_ (.A0(\w[57][22] ),
    .A1(\w[61][22] ),
    .A2(\w[59][22] ),
    .A3(\w[63][22] ),
    .S0(net465),
    .S1(net468),
    .X(_04208_));
 sky130_fd_sc_hd__mux4_2 _14567_ (.A0(_04205_),
    .A1(_04206_),
    .A2(_04207_),
    .A3(_04208_),
    .S0(net458),
    .S1(net455),
    .X(_04209_));
 sky130_fd_sc_hd__mux2i_4 _14568_ (.A0(_04204_),
    .A1(_04209_),
    .S(net542),
    .Y(_12008_));
 sky130_fd_sc_hd__xnor2_1 _14569_ (.A(_02738_),
    .B(_04152_),
    .Y(_12013_));
 sky130_fd_sc_hd__xnor2_1 _14570_ (.A(_03530_),
    .B(_03755_),
    .Y(_04210_));
 sky130_fd_sc_hd__xnor2_2 _14571_ (.A(_03120_),
    .B(_04210_),
    .Y(_12012_));
 sky130_fd_sc_hd__mux4_2 _14572_ (.A0(\w[0][23] ),
    .A1(\w[4][23] ),
    .A2(\w[2][23] ),
    .A3(\w[6][23] ),
    .S0(net386),
    .S1(net393),
    .X(_04211_));
 sky130_fd_sc_hd__mux4_2 _14573_ (.A0(\w[8][23] ),
    .A1(\w[12][23] ),
    .A2(\w[10][23] ),
    .A3(\w[14][23] ),
    .S0(net386),
    .S1(net393),
    .X(_04212_));
 sky130_fd_sc_hd__mux4_2 _14574_ (.A0(\w[16][23] ),
    .A1(\w[20][23] ),
    .A2(\w[18][23] ),
    .A3(\w[22][23] ),
    .S0(net386),
    .S1(net393),
    .X(_04213_));
 sky130_fd_sc_hd__mux4_2 _14575_ (.A0(\w[24][23] ),
    .A1(\w[28][23] ),
    .A2(\w[26][23] ),
    .A3(\w[30][23] ),
    .S0(net386),
    .S1(net393),
    .X(_04214_));
 sky130_fd_sc_hd__mux4_2 _14576_ (.A0(_04211_),
    .A1(_04212_),
    .A2(_04213_),
    .A3(_04214_),
    .S0(net377),
    .S1(net375),
    .X(_04215_));
 sky130_fd_sc_hd__mux4_2 _14577_ (.A0(\w[32][23] ),
    .A1(\w[36][23] ),
    .A2(\w[34][23] ),
    .A3(\w[38][23] ),
    .S0(net384),
    .S1(net391),
    .X(_04216_));
 sky130_fd_sc_hd__mux4_2 _14578_ (.A0(\w[40][23] ),
    .A1(\w[44][23] ),
    .A2(\w[42][23] ),
    .A3(\w[46][23] ),
    .S0(net384),
    .S1(net391),
    .X(_04217_));
 sky130_fd_sc_hd__mux4_2 _14579_ (.A0(\w[48][23] ),
    .A1(\w[52][23] ),
    .A2(\w[50][23] ),
    .A3(\w[54][23] ),
    .S0(net384),
    .S1(net391),
    .X(_04218_));
 sky130_fd_sc_hd__mux4_2 _14580_ (.A0(\w[56][23] ),
    .A1(\w[60][23] ),
    .A2(\w[58][23] ),
    .A3(\w[62][23] ),
    .S0(net384),
    .S1(net391),
    .X(_04219_));
 sky130_fd_sc_hd__mux4_2 _14581_ (.A0(_04216_),
    .A1(_04217_),
    .A2(_04218_),
    .A3(_04219_),
    .S0(net377),
    .S1(net375),
    .X(_04220_));
 sky130_fd_sc_hd__mux2i_4 _14582_ (.A0(_04215_),
    .A1(_04220_),
    .S(net373),
    .Y(_12011_));
 sky130_fd_sc_hd__mux4_2 _14583_ (.A0(\w[1][23] ),
    .A1(\w[5][23] ),
    .A2(\w[3][23] ),
    .A3(\w[7][23] ),
    .S0(net462),
    .S1(net544),
    .X(_04221_));
 sky130_fd_sc_hd__mux4_2 _14584_ (.A0(\w[9][23] ),
    .A1(\w[13][23] ),
    .A2(\w[11][23] ),
    .A3(\w[15][23] ),
    .S0(net462),
    .S1(net544),
    .X(_04222_));
 sky130_fd_sc_hd__mux4_2 _14585_ (.A0(\w[17][23] ),
    .A1(\w[21][23] ),
    .A2(\w[19][23] ),
    .A3(\w[23][23] ),
    .S0(net462),
    .S1(net544),
    .X(_04223_));
 sky130_fd_sc_hd__mux4_2 _14586_ (.A0(\w[25][23] ),
    .A1(\w[29][23] ),
    .A2(\w[27][23] ),
    .A3(\w[31][23] ),
    .S0(net462),
    .S1(net544),
    .X(_04224_));
 sky130_fd_sc_hd__mux4_2 _14587_ (.A0(_04221_),
    .A1(_04222_),
    .A2(_04223_),
    .A3(_04224_),
    .S0(net457),
    .S1(\count16_2[4] ),
    .X(_04225_));
 sky130_fd_sc_hd__mux4_2 _14588_ (.A0(\w[33][23] ),
    .A1(\w[37][23] ),
    .A2(\w[35][23] ),
    .A3(\w[39][23] ),
    .S0(net460),
    .S1(net469),
    .X(_04226_));
 sky130_fd_sc_hd__mux4_2 _14589_ (.A0(\w[41][23] ),
    .A1(\w[45][23] ),
    .A2(\w[43][23] ),
    .A3(\w[47][23] ),
    .S0(net461),
    .S1(net469),
    .X(_04227_));
 sky130_fd_sc_hd__mux4_2 _14590_ (.A0(\w[49][23] ),
    .A1(\w[53][23] ),
    .A2(\w[51][23] ),
    .A3(\w[55][23] ),
    .S0(net461),
    .S1(net469),
    .X(_04228_));
 sky130_fd_sc_hd__mux4_2 _14591_ (.A0(\w[57][23] ),
    .A1(\w[61][23] ),
    .A2(\w[59][23] ),
    .A3(\w[63][23] ),
    .S0(net461),
    .S1(net469),
    .X(_04229_));
 sky130_fd_sc_hd__mux4_2 _14592_ (.A0(_04226_),
    .A1(_04227_),
    .A2(_04228_),
    .A3(_04229_),
    .S0(net457),
    .S1(net543),
    .X(_04230_));
 sky130_fd_sc_hd__mux2i_4 _14593_ (.A0(_04225_),
    .A1(_04230_),
    .S(net453),
    .Y(_12016_));
 sky130_fd_sc_hd__xnor2_1 _14594_ (.A(_02938_),
    .B(_04188_),
    .Y(_12021_));
 sky130_fd_sc_hd__xnor2_1 _14595_ (.A(_03590_),
    .B(_03815_),
    .Y(_04231_));
 sky130_fd_sc_hd__xnor2_1 _14596_ (.A(_03205_),
    .B(_04231_),
    .Y(_12020_));
 sky130_fd_sc_hd__mux4_2 _14597_ (.A0(\w[0][24] ),
    .A1(\w[4][24] ),
    .A2(\w[2][24] ),
    .A3(\w[6][24] ),
    .S0(net381),
    .S1(net389),
    .X(_04232_));
 sky130_fd_sc_hd__mux4_2 _14598_ (.A0(\w[8][24] ),
    .A1(\w[12][24] ),
    .A2(\w[10][24] ),
    .A3(\w[14][24] ),
    .S0(net381),
    .S1(net389),
    .X(_04233_));
 sky130_fd_sc_hd__mux4_2 _14599_ (.A0(\w[16][24] ),
    .A1(\w[20][24] ),
    .A2(\w[18][24] ),
    .A3(\w[22][24] ),
    .S0(net381),
    .S1(net389),
    .X(_04234_));
 sky130_fd_sc_hd__mux4_2 _14600_ (.A0(\w[24][24] ),
    .A1(\w[28][24] ),
    .A2(\w[26][24] ),
    .A3(\w[30][24] ),
    .S0(net381),
    .S1(net389),
    .X(_04235_));
 sky130_fd_sc_hd__mux4_2 _14601_ (.A0(_04232_),
    .A1(_04233_),
    .A2(_04234_),
    .A3(_04235_),
    .S0(net378),
    .S1(net535),
    .X(_04236_));
 sky130_fd_sc_hd__mux4_2 _14602_ (.A0(\w[32][24] ),
    .A1(\w[36][24] ),
    .A2(\w[34][24] ),
    .A3(\w[38][24] ),
    .S0(net382),
    .S1(net389),
    .X(_04237_));
 sky130_fd_sc_hd__mux4_2 _14603_ (.A0(\w[40][24] ),
    .A1(\w[44][24] ),
    .A2(\w[42][24] ),
    .A3(\w[46][24] ),
    .S0(net381),
    .S1(net389),
    .X(_04238_));
 sky130_fd_sc_hd__mux4_2 _14604_ (.A0(\w[48][24] ),
    .A1(\w[52][24] ),
    .A2(\w[50][24] ),
    .A3(\w[54][24] ),
    .S0(net382),
    .S1(net389),
    .X(_04239_));
 sky130_fd_sc_hd__mux4_2 _14605_ (.A0(\w[56][24] ),
    .A1(\w[60][24] ),
    .A2(\w[58][24] ),
    .A3(\w[62][24] ),
    .S0(net382),
    .S1(net389),
    .X(_04240_));
 sky130_fd_sc_hd__mux4_2 _14606_ (.A0(_04237_),
    .A1(_04238_),
    .A2(_04239_),
    .A3(_04240_),
    .S0(net377),
    .S1(net535),
    .X(_04241_));
 sky130_fd_sc_hd__mux2i_4 _14607_ (.A0(_04236_),
    .A1(_04241_),
    .S(net374),
    .Y(_12019_));
 sky130_fd_sc_hd__mux4_2 _14608_ (.A0(\w[1][24] ),
    .A1(\w[5][24] ),
    .A2(\w[3][24] ),
    .A3(\w[7][24] ),
    .S0(net460),
    .S1(net470),
    .X(_04242_));
 sky130_fd_sc_hd__mux4_2 _14609_ (.A0(\w[9][24] ),
    .A1(\w[13][24] ),
    .A2(\w[11][24] ),
    .A3(\w[15][24] ),
    .S0(net460),
    .S1(net470),
    .X(_04243_));
 sky130_fd_sc_hd__mux4_2 _14610_ (.A0(\w[17][24] ),
    .A1(\w[21][24] ),
    .A2(\w[19][24] ),
    .A3(\w[23][24] ),
    .S0(net460),
    .S1(net470),
    .X(_04244_));
 sky130_fd_sc_hd__mux4_2 _14611_ (.A0(\w[25][24] ),
    .A1(\w[29][24] ),
    .A2(\w[27][24] ),
    .A3(\w[31][24] ),
    .S0(net460),
    .S1(net470),
    .X(_04245_));
 sky130_fd_sc_hd__mux4_2 _14612_ (.A0(_04242_),
    .A1(_04243_),
    .A2(_04244_),
    .A3(_04245_),
    .S0(net456),
    .S1(net454),
    .X(_04246_));
 sky130_fd_sc_hd__mux4_2 _14613_ (.A0(\w[33][24] ),
    .A1(\w[37][24] ),
    .A2(\w[35][24] ),
    .A3(\w[39][24] ),
    .S0(net460),
    .S1(net469),
    .X(_04247_));
 sky130_fd_sc_hd__mux4_2 _14614_ (.A0(\w[41][24] ),
    .A1(\w[45][24] ),
    .A2(\w[43][24] ),
    .A3(\w[47][24] ),
    .S0(net460),
    .S1(net469),
    .X(_04248_));
 sky130_fd_sc_hd__mux4_2 _14615_ (.A0(\w[49][24] ),
    .A1(\w[53][24] ),
    .A2(\w[51][24] ),
    .A3(\w[55][24] ),
    .S0(net460),
    .S1(net469),
    .X(_04249_));
 sky130_fd_sc_hd__mux4_2 _14616_ (.A0(\w[57][24] ),
    .A1(\w[61][24] ),
    .A2(\w[59][24] ),
    .A3(\w[63][24] ),
    .S0(net460),
    .S1(net469),
    .X(_04250_));
 sky130_fd_sc_hd__mux4_2 _14617_ (.A0(_04247_),
    .A1(_04248_),
    .A2(_04249_),
    .A3(_04250_),
    .S0(net456),
    .S1(net543),
    .X(_04251_));
 sky130_fd_sc_hd__mux2i_4 _14618_ (.A0(_04246_),
    .A1(_04251_),
    .S(net453),
    .Y(_12024_));
 sky130_fd_sc_hd__xnor2_1 _14619_ (.A(_02738_),
    .B(_03075_),
    .Y(_12029_));
 sky130_fd_sc_hd__xnor2_1 _14620_ (.A(_03645_),
    .B(_03864_),
    .Y(_04252_));
 sky130_fd_sc_hd__xnor2_1 _14621_ (.A(_03275_),
    .B(_04252_),
    .Y(_12028_));
 sky130_fd_sc_hd__mux4_2 _14622_ (.A0(\w[0][25] ),
    .A1(\w[4][25] ),
    .A2(\w[2][25] ),
    .A3(\w[6][25] ),
    .S0(net384),
    .S1(net391),
    .X(_04253_));
 sky130_fd_sc_hd__mux4_2 _14623_ (.A0(\w[8][25] ),
    .A1(\w[12][25] ),
    .A2(\w[10][25] ),
    .A3(\w[14][25] ),
    .S0(net384),
    .S1(net391),
    .X(_04254_));
 sky130_fd_sc_hd__mux4_2 _14624_ (.A0(\w[16][25] ),
    .A1(\w[20][25] ),
    .A2(\w[18][25] ),
    .A3(\w[22][25] ),
    .S0(net384),
    .S1(net391),
    .X(_04255_));
 sky130_fd_sc_hd__mux4_2 _14625_ (.A0(\w[24][25] ),
    .A1(\w[28][25] ),
    .A2(\w[26][25] ),
    .A3(\w[30][25] ),
    .S0(net384),
    .S1(net391),
    .X(_04256_));
 sky130_fd_sc_hd__mux4_2 _14626_ (.A0(_04253_),
    .A1(_04254_),
    .A2(_04255_),
    .A3(_04256_),
    .S0(net377),
    .S1(net375),
    .X(_04257_));
 sky130_fd_sc_hd__mux4_2 _14627_ (.A0(\w[32][25] ),
    .A1(\w[36][25] ),
    .A2(\w[34][25] ),
    .A3(\w[38][25] ),
    .S0(net383),
    .S1(net390),
    .X(_04258_));
 sky130_fd_sc_hd__mux4_2 _14628_ (.A0(\w[40][25] ),
    .A1(\w[44][25] ),
    .A2(\w[42][25] ),
    .A3(\w[46][25] ),
    .S0(net384),
    .S1(net391),
    .X(_04259_));
 sky130_fd_sc_hd__mux4_2 _14629_ (.A0(\w[48][25] ),
    .A1(\w[52][25] ),
    .A2(\w[50][25] ),
    .A3(\w[54][25] ),
    .S0(net384),
    .S1(net391),
    .X(_04260_));
 sky130_fd_sc_hd__mux4_2 _14630_ (.A0(\w[56][25] ),
    .A1(\w[60][25] ),
    .A2(\w[58][25] ),
    .A3(\w[62][25] ),
    .S0(net384),
    .S1(net391),
    .X(_04261_));
 sky130_fd_sc_hd__mux4_2 _14631_ (.A0(_04258_),
    .A1(_04259_),
    .A2(_04260_),
    .A3(_04261_),
    .S0(net377),
    .S1(net375),
    .X(_04262_));
 sky130_fd_sc_hd__mux2i_4 _14632_ (.A0(_04257_),
    .A1(_04262_),
    .S(net373),
    .Y(_12027_));
 sky130_fd_sc_hd__mux4_2 _14633_ (.A0(\w[1][25] ),
    .A1(\w[5][25] ),
    .A2(\w[3][25] ),
    .A3(\w[7][25] ),
    .S0(net465),
    .S1(net468),
    .X(_04263_));
 sky130_fd_sc_hd__mux4_2 _14634_ (.A0(\w[9][25] ),
    .A1(\w[13][25] ),
    .A2(\w[11][25] ),
    .A3(\w[15][25] ),
    .S0(net465),
    .S1(net468),
    .X(_04264_));
 sky130_fd_sc_hd__mux4_2 _14635_ (.A0(\w[17][25] ),
    .A1(\w[21][25] ),
    .A2(\w[19][25] ),
    .A3(\w[23][25] ),
    .S0(net464),
    .S1(net468),
    .X(_04265_));
 sky130_fd_sc_hd__mux4_2 _14636_ (.A0(\w[25][25] ),
    .A1(\w[29][25] ),
    .A2(\w[27][25] ),
    .A3(\w[31][25] ),
    .S0(net464),
    .S1(net468),
    .X(_04266_));
 sky130_fd_sc_hd__mux4_2 _14637_ (.A0(_04263_),
    .A1(_04264_),
    .A2(_04265_),
    .A3(_04266_),
    .S0(net458),
    .S1(net454),
    .X(_04267_));
 sky130_fd_sc_hd__mux4_2 _14638_ (.A0(\w[33][25] ),
    .A1(\w[37][25] ),
    .A2(\w[35][25] ),
    .A3(\w[39][25] ),
    .S0(net464),
    .S1(net468),
    .X(_04268_));
 sky130_fd_sc_hd__mux4_2 _14639_ (.A0(\w[41][25] ),
    .A1(\w[45][25] ),
    .A2(\w[43][25] ),
    .A3(\w[47][25] ),
    .S0(net464),
    .S1(net468),
    .X(_04269_));
 sky130_fd_sc_hd__mux4_2 _14640_ (.A0(\w[49][25] ),
    .A1(\w[53][25] ),
    .A2(\w[51][25] ),
    .A3(\w[55][25] ),
    .S0(net464),
    .S1(net468),
    .X(_04270_));
 sky130_fd_sc_hd__mux4_2 _14641_ (.A0(\w[57][25] ),
    .A1(\w[61][25] ),
    .A2(\w[59][25] ),
    .A3(\w[63][25] ),
    .S0(net464),
    .S1(net468),
    .X(_04271_));
 sky130_fd_sc_hd__mux4_2 _14642_ (.A0(_04268_),
    .A1(_04269_),
    .A2(_04270_),
    .A3(_04271_),
    .S0(\count16_2[3] ),
    .S1(net543),
    .X(_04272_));
 sky130_fd_sc_hd__mux2i_4 _14643_ (.A0(_04267_),
    .A1(_04272_),
    .S(net542),
    .Y(_12032_));
 sky130_fd_sc_hd__xnor2_1 _14644_ (.A(_02938_),
    .B(_03157_),
    .Y(_12037_));
 sky130_fd_sc_hd__xnor2_1 _14645_ (.A(_03709_),
    .B(_03910_),
    .Y(_04273_));
 sky130_fd_sc_hd__xnor2_1 _14646_ (.A(_03344_),
    .B(_04273_),
    .Y(_12036_));
 sky130_fd_sc_hd__mux4_2 _14647_ (.A0(\w[0][26] ),
    .A1(\w[4][26] ),
    .A2(\w[2][26] ),
    .A3(\w[6][26] ),
    .S0(net384),
    .S1(net391),
    .X(_04274_));
 sky130_fd_sc_hd__mux4_2 _14648_ (.A0(\w[8][26] ),
    .A1(\w[12][26] ),
    .A2(\w[10][26] ),
    .A3(\w[14][26] ),
    .S0(net384),
    .S1(net391),
    .X(_04275_));
 sky130_fd_sc_hd__mux4_2 _14649_ (.A0(\w[16][26] ),
    .A1(\w[20][26] ),
    .A2(\w[18][26] ),
    .A3(\w[22][26] ),
    .S0(net384),
    .S1(net391),
    .X(_04276_));
 sky130_fd_sc_hd__mux4_2 _14650_ (.A0(\w[24][26] ),
    .A1(\w[28][26] ),
    .A2(\w[26][26] ),
    .A3(\w[30][26] ),
    .S0(net384),
    .S1(net391),
    .X(_04277_));
 sky130_fd_sc_hd__mux4_2 _14651_ (.A0(_04274_),
    .A1(_04275_),
    .A2(_04276_),
    .A3(_04277_),
    .S0(net377),
    .S1(net375),
    .X(_04278_));
 sky130_fd_sc_hd__mux4_2 _14652_ (.A0(\w[32][26] ),
    .A1(\w[36][26] ),
    .A2(\w[34][26] ),
    .A3(\w[38][26] ),
    .S0(net384),
    .S1(net391),
    .X(_04279_));
 sky130_fd_sc_hd__mux4_2 _14653_ (.A0(\w[40][26] ),
    .A1(\w[44][26] ),
    .A2(\w[42][26] ),
    .A3(\w[46][26] ),
    .S0(net384),
    .S1(net391),
    .X(_04280_));
 sky130_fd_sc_hd__mux4_2 _14654_ (.A0(\w[48][26] ),
    .A1(\w[52][26] ),
    .A2(\w[50][26] ),
    .A3(\w[54][26] ),
    .S0(net384),
    .S1(net391),
    .X(_04281_));
 sky130_fd_sc_hd__mux4_2 _14655_ (.A0(\w[56][26] ),
    .A1(\w[60][26] ),
    .A2(\w[58][26] ),
    .A3(\w[62][26] ),
    .S0(net384),
    .S1(net391),
    .X(_04282_));
 sky130_fd_sc_hd__mux4_2 _14656_ (.A0(_04279_),
    .A1(_04280_),
    .A2(_04281_),
    .A3(_04282_),
    .S0(net377),
    .S1(net375),
    .X(_04283_));
 sky130_fd_sc_hd__mux2i_4 _14657_ (.A0(_04278_),
    .A1(_04283_),
    .S(net373),
    .Y(_12035_));
 sky130_fd_sc_hd__mux4_2 _14658_ (.A0(\w[1][26] ),
    .A1(\w[5][26] ),
    .A2(\w[3][26] ),
    .A3(\w[7][26] ),
    .S0(net462),
    .S1(\count16_2[1] ),
    .X(_04284_));
 sky130_fd_sc_hd__mux4_2 _14659_ (.A0(\w[9][26] ),
    .A1(\w[13][26] ),
    .A2(\w[11][26] ),
    .A3(\w[15][26] ),
    .S0(net462),
    .S1(\count16_2[1] ),
    .X(_04285_));
 sky130_fd_sc_hd__mux4_2 _14660_ (.A0(\w[17][26] ),
    .A1(\w[21][26] ),
    .A2(\w[19][26] ),
    .A3(\w[23][26] ),
    .S0(net462),
    .S1(net544),
    .X(_04286_));
 sky130_fd_sc_hd__mux4_2 _14661_ (.A0(\w[25][26] ),
    .A1(\w[29][26] ),
    .A2(\w[27][26] ),
    .A3(\w[31][26] ),
    .S0(net462),
    .S1(\count16_2[1] ),
    .X(_04287_));
 sky130_fd_sc_hd__mux4_2 _14662_ (.A0(_04284_),
    .A1(_04285_),
    .A2(_04286_),
    .A3(_04287_),
    .S0(net457),
    .S1(\count16_2[4] ),
    .X(_04288_));
 sky130_fd_sc_hd__mux4_2 _14663_ (.A0(\w[33][26] ),
    .A1(\w[37][26] ),
    .A2(\w[35][26] ),
    .A3(\w[39][26] ),
    .S0(net462),
    .S1(net470),
    .X(_04289_));
 sky130_fd_sc_hd__mux4_2 _14664_ (.A0(\w[41][26] ),
    .A1(\w[45][26] ),
    .A2(\w[43][26] ),
    .A3(\w[47][26] ),
    .S0(net462),
    .S1(net470),
    .X(_04290_));
 sky130_fd_sc_hd__mux4_2 _14665_ (.A0(\w[49][26] ),
    .A1(\w[53][26] ),
    .A2(\w[51][26] ),
    .A3(\w[55][26] ),
    .S0(net462),
    .S1(net470),
    .X(_04291_));
 sky130_fd_sc_hd__mux4_2 _14666_ (.A0(\w[57][26] ),
    .A1(\w[61][26] ),
    .A2(\w[59][26] ),
    .A3(\w[63][26] ),
    .S0(net462),
    .S1(net470),
    .X(_04292_));
 sky130_fd_sc_hd__mux4_2 _14667_ (.A0(_04289_),
    .A1(_04290_),
    .A2(_04291_),
    .A3(_04292_),
    .S0(net457),
    .S1(\count16_2[4] ),
    .X(_04293_));
 sky130_fd_sc_hd__mux2i_4 _14668_ (.A0(_04288_),
    .A1(_04293_),
    .S(\count16_2[5] ),
    .Y(_12040_));
 sky130_fd_sc_hd__xnor2_1 _14669_ (.A(_03075_),
    .B(_03239_),
    .Y(_12045_));
 sky130_fd_sc_hd__xnor2_1 _14670_ (.A(_03755_),
    .B(_03956_),
    .Y(_04294_));
 sky130_fd_sc_hd__xnor2_1 _14671_ (.A(_03402_),
    .B(_04294_),
    .Y(_12044_));
 sky130_fd_sc_hd__mux4_2 _14672_ (.A0(\w[0][27] ),
    .A1(\w[4][27] ),
    .A2(\w[2][27] ),
    .A3(\w[6][27] ),
    .S0(net386),
    .S1(net393),
    .X(_04295_));
 sky130_fd_sc_hd__mux4_2 _14673_ (.A0(\w[8][27] ),
    .A1(\w[12][27] ),
    .A2(\w[10][27] ),
    .A3(\w[14][27] ),
    .S0(net386),
    .S1(net393),
    .X(_04296_));
 sky130_fd_sc_hd__mux4_2 _14674_ (.A0(\w[16][27] ),
    .A1(\w[20][27] ),
    .A2(\w[18][27] ),
    .A3(\w[22][27] ),
    .S0(net386),
    .S1(net393),
    .X(_04297_));
 sky130_fd_sc_hd__mux4_2 _14675_ (.A0(\w[24][27] ),
    .A1(\w[28][27] ),
    .A2(\w[26][27] ),
    .A3(\w[30][27] ),
    .S0(net386),
    .S1(net393),
    .X(_04298_));
 sky130_fd_sc_hd__mux4_2 _14676_ (.A0(_04295_),
    .A1(_04296_),
    .A2(_04297_),
    .A3(_04298_),
    .S0(net377),
    .S1(net375),
    .X(_04299_));
 sky130_fd_sc_hd__mux4_2 _14677_ (.A0(\w[32][27] ),
    .A1(\w[36][27] ),
    .A2(\w[34][27] ),
    .A3(\w[38][27] ),
    .S0(net386),
    .S1(net393),
    .X(_04300_));
 sky130_fd_sc_hd__mux4_2 _14678_ (.A0(\w[40][27] ),
    .A1(\w[44][27] ),
    .A2(\w[42][27] ),
    .A3(\w[46][27] ),
    .S0(net386),
    .S1(net393),
    .X(_04301_));
 sky130_fd_sc_hd__mux4_2 _14679_ (.A0(\w[48][27] ),
    .A1(\w[52][27] ),
    .A2(\w[50][27] ),
    .A3(\w[54][27] ),
    .S0(net386),
    .S1(net393),
    .X(_04302_));
 sky130_fd_sc_hd__mux4_2 _14680_ (.A0(\w[56][27] ),
    .A1(\w[60][27] ),
    .A2(\w[58][27] ),
    .A3(\w[62][27] ),
    .S0(net386),
    .S1(net393),
    .X(_04303_));
 sky130_fd_sc_hd__mux4_2 _14681_ (.A0(_04300_),
    .A1(_04301_),
    .A2(_04302_),
    .A3(_04303_),
    .S0(net379),
    .S1(net376),
    .X(_04304_));
 sky130_fd_sc_hd__mux2i_4 _14682_ (.A0(_04299_),
    .A1(_04304_),
    .S(net373),
    .Y(_12043_));
 sky130_fd_sc_hd__mux4_2 _14683_ (.A0(\w[1][27] ),
    .A1(\w[5][27] ),
    .A2(\w[3][27] ),
    .A3(\w[7][27] ),
    .S0(net459),
    .S1(net470),
    .X(_04305_));
 sky130_fd_sc_hd__mux4_2 _14684_ (.A0(\w[9][27] ),
    .A1(\w[13][27] ),
    .A2(\w[11][27] ),
    .A3(\w[15][27] ),
    .S0(net459),
    .S1(net470),
    .X(_04306_));
 sky130_fd_sc_hd__mux4_2 _14685_ (.A0(\w[17][27] ),
    .A1(\w[21][27] ),
    .A2(\w[19][27] ),
    .A3(\w[23][27] ),
    .S0(net459),
    .S1(net470),
    .X(_04307_));
 sky130_fd_sc_hd__mux4_2 _14686_ (.A0(\w[25][27] ),
    .A1(\w[29][27] ),
    .A2(\w[27][27] ),
    .A3(\w[31][27] ),
    .S0(net459),
    .S1(net470),
    .X(_04308_));
 sky130_fd_sc_hd__mux4_2 _14687_ (.A0(_04305_),
    .A1(_04306_),
    .A2(_04307_),
    .A3(_04308_),
    .S0(net456),
    .S1(net454),
    .X(_04309_));
 sky130_fd_sc_hd__mux4_2 _14688_ (.A0(\w[33][27] ),
    .A1(\w[37][27] ),
    .A2(\w[35][27] ),
    .A3(\w[39][27] ),
    .S0(net460),
    .S1(net469),
    .X(_04310_));
 sky130_fd_sc_hd__mux4_2 _14689_ (.A0(\w[41][27] ),
    .A1(\w[45][27] ),
    .A2(\w[43][27] ),
    .A3(\w[47][27] ),
    .S0(net460),
    .S1(net469),
    .X(_04311_));
 sky130_fd_sc_hd__mux4_2 _14690_ (.A0(\w[49][27] ),
    .A1(\w[53][27] ),
    .A2(\w[51][27] ),
    .A3(\w[55][27] ),
    .S0(net460),
    .S1(net469),
    .X(_04312_));
 sky130_fd_sc_hd__mux4_2 _14691_ (.A0(\w[57][27] ),
    .A1(\w[61][27] ),
    .A2(\w[59][27] ),
    .A3(\w[63][27] ),
    .S0(net460),
    .S1(net469),
    .X(_04313_));
 sky130_fd_sc_hd__mux4_2 _14692_ (.A0(_04310_),
    .A1(_04311_),
    .A2(_04312_),
    .A3(_04313_),
    .S0(net456),
    .S1(net454),
    .X(_04314_));
 sky130_fd_sc_hd__mux2i_4 _14693_ (.A0(_04309_),
    .A1(_04314_),
    .S(net453),
    .Y(_12048_));
 sky130_fd_sc_hd__xnor2_1 _14694_ (.A(_03157_),
    .B(_03309_),
    .Y(_12053_));
 sky130_fd_sc_hd__xnor2_1 _14695_ (.A(_03460_),
    .B(_03815_),
    .Y(_04315_));
 sky130_fd_sc_hd__xnor2_1 _14696_ (.A(_02824_),
    .B(_04315_),
    .Y(_12052_));
 sky130_fd_sc_hd__mux4_2 _14697_ (.A0(\w[0][28] ),
    .A1(\w[4][28] ),
    .A2(\w[2][28] ),
    .A3(\w[6][28] ),
    .S0(net386),
    .S1(net393),
    .X(_04316_));
 sky130_fd_sc_hd__mux4_2 _14698_ (.A0(\w[8][28] ),
    .A1(\w[12][28] ),
    .A2(\w[10][28] ),
    .A3(\w[14][28] ),
    .S0(net386),
    .S1(net393),
    .X(_04317_));
 sky130_fd_sc_hd__mux4_2 _14699_ (.A0(\w[16][28] ),
    .A1(\w[20][28] ),
    .A2(\w[18][28] ),
    .A3(\w[22][28] ),
    .S0(net386),
    .S1(net393),
    .X(_04318_));
 sky130_fd_sc_hd__mux4_2 _14700_ (.A0(\w[24][28] ),
    .A1(\w[28][28] ),
    .A2(\w[26][28] ),
    .A3(\w[30][28] ),
    .S0(net386),
    .S1(net393),
    .X(_04319_));
 sky130_fd_sc_hd__mux4_2 _14701_ (.A0(_04316_),
    .A1(_04317_),
    .A2(_04318_),
    .A3(_04319_),
    .S0(net377),
    .S1(net375),
    .X(_04320_));
 sky130_fd_sc_hd__mux4_2 _14702_ (.A0(\w[32][28] ),
    .A1(\w[36][28] ),
    .A2(\w[34][28] ),
    .A3(\w[38][28] ),
    .S0(net384),
    .S1(net391),
    .X(_04321_));
 sky130_fd_sc_hd__mux4_2 _14703_ (.A0(\w[40][28] ),
    .A1(\w[44][28] ),
    .A2(\w[42][28] ),
    .A3(\w[46][28] ),
    .S0(net384),
    .S1(net391),
    .X(_04322_));
 sky130_fd_sc_hd__mux4_2 _14704_ (.A0(\w[48][28] ),
    .A1(\w[52][28] ),
    .A2(\w[50][28] ),
    .A3(\w[54][28] ),
    .S0(net384),
    .S1(net391),
    .X(_04323_));
 sky130_fd_sc_hd__mux4_2 _14705_ (.A0(\w[56][28] ),
    .A1(\w[60][28] ),
    .A2(\w[58][28] ),
    .A3(\w[62][28] ),
    .S0(net384),
    .S1(net391),
    .X(_04324_));
 sky130_fd_sc_hd__mux4_2 _14706_ (.A0(_04321_),
    .A1(_04322_),
    .A2(_04323_),
    .A3(_04324_),
    .S0(net377),
    .S1(net375),
    .X(_04325_));
 sky130_fd_sc_hd__mux2i_4 _14707_ (.A0(_04320_),
    .A1(_04325_),
    .S(net373),
    .Y(_12051_));
 sky130_fd_sc_hd__mux4_2 _14708_ (.A0(\w[1][28] ),
    .A1(\w[5][28] ),
    .A2(\w[3][28] ),
    .A3(\w[7][28] ),
    .S0(net462),
    .S1(net544),
    .X(_04326_));
 sky130_fd_sc_hd__mux4_2 _14709_ (.A0(\w[9][28] ),
    .A1(\w[13][28] ),
    .A2(\w[11][28] ),
    .A3(\w[15][28] ),
    .S0(net462),
    .S1(net544),
    .X(_04327_));
 sky130_fd_sc_hd__mux4_2 _14710_ (.A0(\w[17][28] ),
    .A1(\w[21][28] ),
    .A2(\w[19][28] ),
    .A3(\w[23][28] ),
    .S0(net462),
    .S1(net544),
    .X(_04328_));
 sky130_fd_sc_hd__mux4_2 _14711_ (.A0(\w[25][28] ),
    .A1(\w[29][28] ),
    .A2(\w[27][28] ),
    .A3(\w[31][28] ),
    .S0(net462),
    .S1(net544),
    .X(_04329_));
 sky130_fd_sc_hd__mux4_2 _14712_ (.A0(_04326_),
    .A1(_04327_),
    .A2(_04328_),
    .A3(_04329_),
    .S0(net457),
    .S1(\count16_2[4] ),
    .X(_04330_));
 sky130_fd_sc_hd__mux4_2 _14713_ (.A0(\w[33][28] ),
    .A1(\w[37][28] ),
    .A2(\w[35][28] ),
    .A3(\w[39][28] ),
    .S0(net462),
    .S1(net471),
    .X(_04331_));
 sky130_fd_sc_hd__mux4_2 _14714_ (.A0(\w[41][28] ),
    .A1(\w[45][28] ),
    .A2(\w[43][28] ),
    .A3(\w[47][28] ),
    .S0(net462),
    .S1(net471),
    .X(_04332_));
 sky130_fd_sc_hd__mux4_2 _14715_ (.A0(\w[49][28] ),
    .A1(\w[53][28] ),
    .A2(\w[51][28] ),
    .A3(\w[55][28] ),
    .S0(net462),
    .S1(net471),
    .X(_04333_));
 sky130_fd_sc_hd__mux4_2 _14716_ (.A0(\w[57][28] ),
    .A1(\w[61][28] ),
    .A2(\w[59][28] ),
    .A3(\w[63][28] ),
    .S0(net462),
    .S1(net471),
    .X(_04334_));
 sky130_fd_sc_hd__mux4_2 _14717_ (.A0(_04331_),
    .A1(_04332_),
    .A2(_04333_),
    .A3(_04334_),
    .S0(net457),
    .S1(\count16_2[4] ),
    .X(_04335_));
 sky130_fd_sc_hd__mux2i_4 _14718_ (.A0(_04330_),
    .A1(_04335_),
    .S(net453),
    .Y(_12056_));
 sky130_fd_sc_hd__xnor2_1 _14719_ (.A(_03239_),
    .B(_03378_),
    .Y(_12061_));
 sky130_fd_sc_hd__xnor2_1 _14720_ (.A(_02976_),
    .B(_03519_),
    .Y(_12060_));
 sky130_fd_sc_hd__mux4_2 _14721_ (.A0(\w[0][29] ),
    .A1(\w[4][29] ),
    .A2(\w[2][29] ),
    .A3(\w[6][29] ),
    .S0(net380),
    .S1(net388),
    .X(_04336_));
 sky130_fd_sc_hd__mux4_2 _14722_ (.A0(\w[8][29] ),
    .A1(\w[12][29] ),
    .A2(\w[10][29] ),
    .A3(\w[14][29] ),
    .S0(net380),
    .S1(net388),
    .X(_04337_));
 sky130_fd_sc_hd__mux4_2 _14723_ (.A0(\w[16][29] ),
    .A1(\w[20][29] ),
    .A2(\w[18][29] ),
    .A3(\w[22][29] ),
    .S0(net380),
    .S1(net388),
    .X(_04338_));
 sky130_fd_sc_hd__mux4_2 _14724_ (.A0(\w[24][29] ),
    .A1(\w[28][29] ),
    .A2(\w[26][29] ),
    .A3(\w[30][29] ),
    .S0(net380),
    .S1(net388),
    .X(_04339_));
 sky130_fd_sc_hd__mux4_2 _14725_ (.A0(_04336_),
    .A1(_04337_),
    .A2(_04338_),
    .A3(_04339_),
    .S0(net379),
    .S1(net376),
    .X(_04340_));
 sky130_fd_sc_hd__mux4_2 _14726_ (.A0(\w[32][29] ),
    .A1(\w[36][29] ),
    .A2(\w[34][29] ),
    .A3(\w[38][29] ),
    .S0(net380),
    .S1(net388),
    .X(_04341_));
 sky130_fd_sc_hd__mux4_2 _14727_ (.A0(\w[40][29] ),
    .A1(\w[44][29] ),
    .A2(\w[42][29] ),
    .A3(\w[46][29] ),
    .S0(net380),
    .S1(net388),
    .X(_04342_));
 sky130_fd_sc_hd__mux4_2 _14728_ (.A0(\w[48][29] ),
    .A1(\w[52][29] ),
    .A2(\w[50][29] ),
    .A3(\w[54][29] ),
    .S0(net380),
    .S1(net388),
    .X(_04343_));
 sky130_fd_sc_hd__mux4_2 _14729_ (.A0(\w[56][29] ),
    .A1(\w[60][29] ),
    .A2(\w[58][29] ),
    .A3(\w[62][29] ),
    .S0(net380),
    .S1(net388),
    .X(_04344_));
 sky130_fd_sc_hd__mux4_2 _14730_ (.A0(_04341_),
    .A1(_04342_),
    .A2(_04343_),
    .A3(_04344_),
    .S0(net379),
    .S1(net376),
    .X(_04345_));
 sky130_fd_sc_hd__mux2i_4 _14731_ (.A0(_04340_),
    .A1(_04345_),
    .S(net373),
    .Y(_12059_));
 sky130_fd_sc_hd__mux4_2 _14732_ (.A0(\w[1][29] ),
    .A1(\w[5][29] ),
    .A2(\w[3][29] ),
    .A3(\w[7][29] ),
    .S0(net466),
    .S1(\count16_2[1] ),
    .X(_04346_));
 sky130_fd_sc_hd__mux4_2 _14733_ (.A0(\w[9][29] ),
    .A1(\w[13][29] ),
    .A2(\w[11][29] ),
    .A3(\w[15][29] ),
    .S0(net466),
    .S1(\count16_2[1] ),
    .X(_04347_));
 sky130_fd_sc_hd__mux4_2 _14734_ (.A0(\w[17][29] ),
    .A1(\w[21][29] ),
    .A2(\w[19][29] ),
    .A3(\w[23][29] ),
    .S0(net466),
    .S1(\count16_2[1] ),
    .X(_04348_));
 sky130_fd_sc_hd__mux4_2 _14735_ (.A0(\w[25][29] ),
    .A1(\w[29][29] ),
    .A2(\w[27][29] ),
    .A3(\w[31][29] ),
    .S0(net466),
    .S1(\count16_2[1] ),
    .X(_04349_));
 sky130_fd_sc_hd__mux4_2 _14736_ (.A0(_04346_),
    .A1(_04347_),
    .A2(_04348_),
    .A3(_04349_),
    .S0(net457),
    .S1(\count16_2[4] ),
    .X(_04350_));
 sky130_fd_sc_hd__mux4_2 _14737_ (.A0(\w[33][29] ),
    .A1(\w[37][29] ),
    .A2(\w[35][29] ),
    .A3(\w[39][29] ),
    .S0(net466),
    .S1(net471),
    .X(_04351_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1427 ();
 sky130_fd_sc_hd__mux4_2 _14739_ (.A0(\w[41][29] ),
    .A1(\w[45][29] ),
    .A2(\w[43][29] ),
    .A3(\w[47][29] ),
    .S0(net466),
    .S1(net471),
    .X(_04353_));
 sky130_fd_sc_hd__mux4_2 _14740_ (.A0(\w[49][29] ),
    .A1(\w[53][29] ),
    .A2(\w[51][29] ),
    .A3(\w[55][29] ),
    .S0(net466),
    .S1(net471),
    .X(_04354_));
 sky130_fd_sc_hd__mux4_2 _14741_ (.A0(\w[57][29] ),
    .A1(\w[61][29] ),
    .A2(\w[59][29] ),
    .A3(\w[63][29] ),
    .S0(net466),
    .S1(net471),
    .X(_04355_));
 sky130_fd_sc_hd__mux4_2 _14742_ (.A0(_04351_),
    .A1(_04353_),
    .A2(_04354_),
    .A3(_04355_),
    .S0(net457),
    .S1(\count16_2[4] ),
    .X(_04356_));
 sky130_fd_sc_hd__mux2i_1 _14743_ (.A0(_04350_),
    .A1(_04356_),
    .S(\count16_2[5] ),
    .Y(_12064_));
 sky130_fd_sc_hd__xnor2_1 _14744_ (.A(_02788_),
    .B(_03309_),
    .Y(_12069_));
 sky130_fd_sc_hd__xnor2_1 _14745_ (.A(_03098_),
    .B(_03579_),
    .Y(_12068_));
 sky130_fd_sc_hd__mux4_2 _14746_ (.A0(\w[0][30] ),
    .A1(\w[4][30] ),
    .A2(\w[2][30] ),
    .A3(\w[6][30] ),
    .S0(net380),
    .S1(net388),
    .X(_04357_));
 sky130_fd_sc_hd__mux4_2 _14747_ (.A0(\w[8][30] ),
    .A1(\w[12][30] ),
    .A2(\w[10][30] ),
    .A3(\w[14][30] ),
    .S0(net380),
    .S1(net388),
    .X(_04358_));
 sky130_fd_sc_hd__mux4_2 _14748_ (.A0(\w[16][30] ),
    .A1(\w[20][30] ),
    .A2(\w[18][30] ),
    .A3(\w[22][30] ),
    .S0(net380),
    .S1(net388),
    .X(_04359_));
 sky130_fd_sc_hd__mux4_2 _14749_ (.A0(\w[24][30] ),
    .A1(\w[28][30] ),
    .A2(\w[26][30] ),
    .A3(\w[30][30] ),
    .S0(net380),
    .S1(net388),
    .X(_04360_));
 sky130_fd_sc_hd__mux4_2 _14750_ (.A0(_04357_),
    .A1(_04358_),
    .A2(_04359_),
    .A3(_04360_),
    .S0(net379),
    .S1(net376),
    .X(_04361_));
 sky130_fd_sc_hd__mux4_2 _14751_ (.A0(\w[32][30] ),
    .A1(\w[36][30] ),
    .A2(\w[34][30] ),
    .A3(\w[38][30] ),
    .S0(net380),
    .S1(net388),
    .X(_04362_));
 sky130_fd_sc_hd__mux4_2 _14752_ (.A0(\w[40][30] ),
    .A1(\w[44][30] ),
    .A2(\w[42][30] ),
    .A3(\w[46][30] ),
    .S0(net380),
    .S1(net388),
    .X(_04363_));
 sky130_fd_sc_hd__mux4_2 _14753_ (.A0(\w[48][30] ),
    .A1(\w[52][30] ),
    .A2(\w[50][30] ),
    .A3(\w[54][30] ),
    .S0(net380),
    .S1(net388),
    .X(_04364_));
 sky130_fd_sc_hd__mux4_2 _14754_ (.A0(\w[56][30] ),
    .A1(\w[60][30] ),
    .A2(\w[58][30] ),
    .A3(\w[62][30] ),
    .S0(net380),
    .S1(net388),
    .X(_04365_));
 sky130_fd_sc_hd__mux4_2 _14755_ (.A0(_04362_),
    .A1(_04363_),
    .A2(_04364_),
    .A3(_04365_),
    .S0(net379),
    .S1(net376),
    .X(_04366_));
 sky130_fd_sc_hd__mux2i_4 _14756_ (.A0(_04361_),
    .A1(_04366_),
    .S(net373),
    .Y(_12067_));
 sky130_fd_sc_hd__mux4_2 _14757_ (.A0(\w[1][30] ),
    .A1(\w[5][30] ),
    .A2(\w[3][30] ),
    .A3(\w[7][30] ),
    .S0(net466),
    .S1(net471),
    .X(_04367_));
 sky130_fd_sc_hd__mux4_2 _14758_ (.A0(\w[9][30] ),
    .A1(\w[13][30] ),
    .A2(\w[11][30] ),
    .A3(\w[15][30] ),
    .S0(net466),
    .S1(net471),
    .X(_04368_));
 sky130_fd_sc_hd__mux4_2 _14759_ (.A0(\w[17][30] ),
    .A1(\w[21][30] ),
    .A2(\w[19][30] ),
    .A3(\w[23][30] ),
    .S0(net466),
    .S1(net471),
    .X(_04369_));
 sky130_fd_sc_hd__mux4_2 _14760_ (.A0(\w[25][30] ),
    .A1(\w[29][30] ),
    .A2(\w[27][30] ),
    .A3(\w[31][30] ),
    .S0(net466),
    .S1(net471),
    .X(_04370_));
 sky130_fd_sc_hd__mux4_2 _14761_ (.A0(_04367_),
    .A1(_04368_),
    .A2(_04369_),
    .A3(_04370_),
    .S0(net457),
    .S1(\count16_2[4] ),
    .X(_04371_));
 sky130_fd_sc_hd__mux4_2 _14762_ (.A0(\w[33][30] ),
    .A1(\w[37][30] ),
    .A2(\w[35][30] ),
    .A3(\w[39][30] ),
    .S0(net466),
    .S1(net471),
    .X(_04372_));
 sky130_fd_sc_hd__mux4_2 _14763_ (.A0(\w[41][30] ),
    .A1(\w[45][30] ),
    .A2(\w[43][30] ),
    .A3(\w[47][30] ),
    .S0(net466),
    .S1(net471),
    .X(_04373_));
 sky130_fd_sc_hd__mux4_2 _14764_ (.A0(\w[49][30] ),
    .A1(\w[53][30] ),
    .A2(\w[51][30] ),
    .A3(\w[55][30] ),
    .S0(net466),
    .S1(net471),
    .X(_04374_));
 sky130_fd_sc_hd__mux4_2 _14765_ (.A0(\w[57][30] ),
    .A1(\w[61][30] ),
    .A2(\w[59][30] ),
    .A3(\w[63][30] ),
    .S0(net466),
    .S1(net471),
    .X(_04375_));
 sky130_fd_sc_hd__mux4_2 _14766_ (.A0(_04372_),
    .A1(_04373_),
    .A2(_04374_),
    .A3(_04375_),
    .S0(net457),
    .S1(net455),
    .X(_04376_));
 sky130_fd_sc_hd__mux2i_1 _14767_ (.A0(_04371_),
    .A1(_04376_),
    .S(\count16_2[5] ),
    .Y(_12072_));
 sky130_fd_sc_hd__a21o_1 _14768_ (.A1(\hash.CA2.a_dash[0] ),
    .A2(_12922_),
    .B1(\hash.CA2.b_dash[0] ),
    .X(_04377_));
 sky130_fd_sc_hd__o21ai_1 _14769_ (.A1(\hash.CA2.a_dash[0] ),
    .A2(_12922_),
    .B1(_04377_),
    .Y(_12077_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1424 ();
 sky130_fd_sc_hd__xnor2_4 _14773_ (.A(\hash.CA2.S1.X[6] ),
    .B(\hash.CA2.S1.X[25] ),
    .Y(_04381_));
 sky130_fd_sc_hd__xnor2_2 _14774_ (.A(_04381_),
    .B(\hash.CA2.S1.X[11] ),
    .Y(_13230_));
 sky130_fd_sc_hd__a21o_1 _14775_ (.A1(_12956_),
    .A2(_12953_),
    .B1(_12955_),
    .X(_04382_));
 sky130_fd_sc_hd__a21oi_1 _14776_ (.A1(_12958_),
    .A2(_04382_),
    .B1(_12957_),
    .Y(_04383_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1423 ();
 sky130_fd_sc_hd__nand2_1 _14778_ (.A(_12962_),
    .B(_12964_),
    .Y(_04385_));
 sky130_fd_sc_hd__nand2_1 _14779_ (.A(_12962_),
    .B(_12963_),
    .Y(_04386_));
 sky130_fd_sc_hd__o21ai_0 _14780_ (.A1(_04383_),
    .A2(_04385_),
    .B1(_04386_),
    .Y(_04387_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1422 ();
 sky130_fd_sc_hd__nand3_1 _14782_ (.A(_12946_),
    .B(_12950_),
    .C(_12952_),
    .Y(_04389_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1421 ();
 sky130_fd_sc_hd__nor2_1 _14784_ (.A(_12948_),
    .B(_12947_),
    .Y(_04391_));
 sky130_fd_sc_hd__a21o_1 _14785_ (.A1(_12952_),
    .A2(_12945_),
    .B1(_12951_),
    .X(_04392_));
 sky130_fd_sc_hd__a21oi_2 _14786_ (.A1(_12950_),
    .A2(_04392_),
    .B1(_12949_),
    .Y(_04393_));
 sky130_fd_sc_hd__o21a_4 _14787_ (.A1(_04389_),
    .A2(_04391_),
    .B1(_04393_),
    .X(_04394_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1420 ();
 sky130_fd_sc_hd__or2_4 _14789_ (.A(_12930_),
    .B(_12929_),
    .X(_04396_));
 sky130_fd_sc_hd__a21o_4 _14790_ (.A1(_12928_),
    .A2(_04396_),
    .B1(_12927_),
    .X(_04397_));
 sky130_fd_sc_hd__a211oi_4 _14791_ (.A1(_12924_),
    .A2(_12081_),
    .B1(_12923_),
    .C1(_12935_),
    .Y(_04398_));
 sky130_fd_sc_hd__o211ai_1 _14792_ (.A1(_12936_),
    .A2(_12935_),
    .B1(_12932_),
    .C1(_12934_),
    .Y(_04399_));
 sky130_fd_sc_hd__a21oi_2 _14793_ (.A1(_12932_),
    .A2(_12933_),
    .B1(_12931_),
    .Y(_04400_));
 sky130_fd_sc_hd__nor2_1 _14794_ (.A(_12927_),
    .B(_12929_),
    .Y(_04401_));
 sky130_fd_sc_hd__o211ai_1 _14795_ (.A1(_04398_),
    .A2(_04399_),
    .B1(_04400_),
    .C1(_04401_),
    .Y(_04402_));
 sky130_fd_sc_hd__clkinv_1 _14796_ (.A(_12944_),
    .Y(_04403_));
 sky130_fd_sc_hd__nand2_4 _14797_ (.A(_12938_),
    .B(_12942_),
    .Y(_04404_));
 sky130_fd_sc_hd__nor2_1 _14798_ (.A(_04403_),
    .B(_04404_),
    .Y(_04405_));
 sky130_fd_sc_hd__and4_4 _14799_ (.A(_12940_),
    .B(_04397_),
    .C(_04402_),
    .D(_04405_),
    .X(_04406_));
 sky130_fd_sc_hd__nand2_2 _14800_ (.A(_12944_),
    .B(_12939_),
    .Y(_04407_));
 sky130_fd_sc_hd__a21oi_4 _14801_ (.A1(_12942_),
    .A2(_12937_),
    .B1(_12941_),
    .Y(_04408_));
 sky130_fd_sc_hd__o22ai_4 _14802_ (.A1(_04404_),
    .A2(_04407_),
    .B1(_04408_),
    .B2(_04403_),
    .Y(_04409_));
 sky130_fd_sc_hd__nor2_1 _14803_ (.A(_12943_),
    .B(_04409_),
    .Y(_04410_));
 sky130_fd_sc_hd__nor4bb_4 _14804_ (.A(_12947_),
    .B(_04406_),
    .C_N(_04410_),
    .D_N(_04393_),
    .Y(_04411_));
 sky130_fd_sc_hd__nand3_1 _14805_ (.A(_12954_),
    .B(_12956_),
    .C(_12958_),
    .Y(_04412_));
 sky130_fd_sc_hd__or4_4 _14806_ (.A(_04411_),
    .B(_04385_),
    .C(_04412_),
    .D(_04394_),
    .X(_04413_));
 sky130_fd_sc_hd__nand2b_1 _14807_ (.A_N(_04387_),
    .B(_04413_),
    .Y(_04414_));
 sky130_fd_sc_hd__o21ai_2 _14808_ (.A1(_12961_),
    .A2(_04414_),
    .B1(_12960_),
    .Y(_04415_));
 sky130_fd_sc_hd__nor2_2 _14809_ (.A(_12966_),
    .B(_12959_),
    .Y(_04416_));
 sky130_fd_sc_hd__nor3_1 _14810_ (.A(_12959_),
    .B(_12961_),
    .C(_04387_),
    .Y(_04417_));
 sky130_fd_sc_hd__o21ai_0 _14811_ (.A1(_12960_),
    .A2(_12959_),
    .B1(_12966_),
    .Y(_04418_));
 sky130_fd_sc_hd__a21oi_4 _14812_ (.A1(_04413_),
    .A2(_04417_),
    .B1(_04418_),
    .Y(_04419_));
 sky130_fd_sc_hd__a21oi_4 _14813_ (.A1(_04415_),
    .A2(_04416_),
    .B1(_04419_),
    .Y(_04420_));
 sky130_fd_sc_hd__xor2_4 _14814_ (.A(_12924_),
    .B(_12081_),
    .X(_04421_));
 sky130_fd_sc_hd__o31a_1 _14815_ (.A1(_12932_),
    .A2(_12929_),
    .A3(_12931_),
    .B1(_04396_),
    .X(_04422_));
 sky130_fd_sc_hd__a211oi_2 _14816_ (.A1(_12080_),
    .A2(_12926_),
    .B1(_12923_),
    .C1(_12925_),
    .Y(_04423_));
 sky130_fd_sc_hd__o211ai_1 _14817_ (.A1(_12924_),
    .A2(_12923_),
    .B1(_12936_),
    .C1(_12934_),
    .Y(_04424_));
 sky130_fd_sc_hd__a21oi_1 _14818_ (.A1(_12934_),
    .A2(_12935_),
    .B1(_12933_),
    .Y(_04425_));
 sky130_fd_sc_hd__nor2_1 _14819_ (.A(_12929_),
    .B(_12931_),
    .Y(_04426_));
 sky130_fd_sc_hd__o211ai_1 _14820_ (.A1(_04424_),
    .A2(_04423_),
    .B1(_04425_),
    .C1(_04426_),
    .Y(_04427_));
 sky130_fd_sc_hd__nand2_4 _14821_ (.A(_04422_),
    .B(_04427_),
    .Y(_04428_));
 sky130_fd_sc_hd__nand2_1 _14822_ (.A(_12928_),
    .B(_12940_),
    .Y(_04429_));
 sky130_fd_sc_hd__nor2_1 _14823_ (.A(_04404_),
    .B(_04429_),
    .Y(_04430_));
 sky130_fd_sc_hd__nand2_1 _14824_ (.A(_12944_),
    .B(_04430_),
    .Y(_04431_));
 sky130_fd_sc_hd__a21oi_2 _14825_ (.A1(_12940_),
    .A2(_12927_),
    .B1(_12939_),
    .Y(_04432_));
 sky130_fd_sc_hd__o21ai_4 _14826_ (.A1(_04404_),
    .A2(_04432_),
    .B1(_04408_),
    .Y(_04433_));
 sky130_fd_sc_hd__a21oi_1 _14827_ (.A1(_12944_),
    .A2(_04433_),
    .B1(_12943_),
    .Y(_04434_));
 sky130_fd_sc_hd__o21ai_2 _14828_ (.A1(_04428_),
    .A2(_04431_),
    .B1(_04434_),
    .Y(_04435_));
 sky130_fd_sc_hd__a21oi_4 _14829_ (.A1(_12948_),
    .A2(_04435_),
    .B1(_12947_),
    .Y(_04436_));
 sky130_fd_sc_hd__xnor2_4 _14830_ (.A(_12946_),
    .B(_04436_),
    .Y(_04437_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1419 ();
 sky130_fd_sc_hd__xor2_1 _14832_ (.A(_04421_),
    .B(_04437_),
    .X(_04439_));
 sky130_fd_sc_hd__xnor2_2 _14833_ (.A(_04420_),
    .B(_04439_),
    .Y(_12075_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1418 ();
 sky130_fd_sc_hd__nor2_4 _14835_ (.A(net340),
    .B(_13235_),
    .Y(_00658_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1417 ();
 sky130_fd_sc_hd__a21o_1 _14837_ (.A1(\hash.CA2.a_dash[1] ),
    .A2(_12082_),
    .B1(\hash.CA2.b_dash[1] ),
    .X(_04442_));
 sky130_fd_sc_hd__o21ai_0 _14838_ (.A1(\hash.CA2.a_dash[1] ),
    .A2(_12082_),
    .B1(_04442_),
    .Y(_12089_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1414 ();
 sky130_fd_sc_hd__xnor2_4 _14842_ (.A(\hash.CA2.S1.X[7] ),
    .B(\hash.CA2.S1.X[26] ),
    .Y(_04446_));
 sky130_fd_sc_hd__xnor2_4 _14843_ (.A(\hash.CA2.S1.X[12] ),
    .B(_04446_),
    .Y(_13237_));
 sky130_fd_sc_hd__inv_2 _14844_ (.A(net1089),
    .Y(_12085_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1413 ();
 sky130_fd_sc_hd__mux2_2 _14846_ (.A0(\hash.CA2.f_dash[1] ),
    .A1(\hash.CA2.e_dash[1] ),
    .S(\hash.CA2.S1.X[1] ),
    .X(_13236_));
 sky130_fd_sc_hd__inv_1 _14847_ (.A(_13236_),
    .Y(_12084_));
 sky130_fd_sc_hd__a21o_1 _14848_ (.A1(_12954_),
    .A2(_12949_),
    .B1(_12953_),
    .X(_04448_));
 sky130_fd_sc_hd__a21o_1 _14849_ (.A1(_12956_),
    .A2(_04448_),
    .B1(_12955_),
    .X(_04449_));
 sky130_fd_sc_hd__a21o_1 _14850_ (.A1(_12958_),
    .A2(_04449_),
    .B1(_12957_),
    .X(_04450_));
 sky130_fd_sc_hd__a21o_1 _14851_ (.A1(_12948_),
    .A2(_12943_),
    .B1(_12947_),
    .X(_04451_));
 sky130_fd_sc_hd__a21o_1 _14852_ (.A1(_12946_),
    .A2(_04451_),
    .B1(_12945_),
    .X(_04452_));
 sky130_fd_sc_hd__a21o_4 _14853_ (.A1(_12952_),
    .A2(_04452_),
    .B1(_12951_),
    .X(_04453_));
 sky130_fd_sc_hd__inv_1 _14854_ (.A(_12964_),
    .Y(_04454_));
 sky130_fd_sc_hd__nand4_1 _14855_ (.A(_12950_),
    .B(_12954_),
    .C(_12956_),
    .D(_12958_),
    .Y(_04455_));
 sky130_fd_sc_hd__nor2_2 _14856_ (.A(_04454_),
    .B(_04455_),
    .Y(_04456_));
 sky130_fd_sc_hd__a22oi_1 _14857_ (.A1(_12964_),
    .A2(_04450_),
    .B1(_04453_),
    .B2(_04456_),
    .Y(_04457_));
 sky130_fd_sc_hd__and3_4 _14858_ (.A(_04422_),
    .B(_04427_),
    .C(_04430_),
    .X(_04458_));
 sky130_fd_sc_hd__nand4_1 _14859_ (.A(_12946_),
    .B(_12944_),
    .C(_12948_),
    .D(_12952_),
    .Y(_04459_));
 sky130_fd_sc_hd__inv_1 _14860_ (.A(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__o211ai_1 _14861_ (.A1(_04433_),
    .A2(_04458_),
    .B1(_04460_),
    .C1(_04456_),
    .Y(_04461_));
 sky130_fd_sc_hd__nor3_1 _14862_ (.A(_12959_),
    .B(_12961_),
    .C(_12963_),
    .Y(_04462_));
 sky130_fd_sc_hd__nand3_2 _14863_ (.A(_04457_),
    .B(_04461_),
    .C(_04462_),
    .Y(_04463_));
 sky130_fd_sc_hd__o21ai_0 _14864_ (.A1(_12962_),
    .A2(_12961_),
    .B1(_12960_),
    .Y(_04464_));
 sky130_fd_sc_hd__nand2b_2 _14865_ (.A_N(_12959_),
    .B(_04464_),
    .Y(_04465_));
 sky130_fd_sc_hd__a31oi_2 _14866_ (.A1(_12966_),
    .A2(_04463_),
    .A3(_04465_),
    .B1(_12965_),
    .Y(_04466_));
 sky130_fd_sc_hd__xnor2_4 _14867_ (.A(_12970_),
    .B(_04466_),
    .Y(_04467_));
 sky130_fd_sc_hd__a21o_1 _14868_ (.A1(_12080_),
    .A2(_12926_),
    .B1(_12925_),
    .X(_04468_));
 sky130_fd_sc_hd__a21oi_2 _14869_ (.A1(_12924_),
    .A2(_04468_),
    .B1(_12923_),
    .Y(_04469_));
 sky130_fd_sc_hd__xnor2_4 _14870_ (.A(_12936_),
    .B(_04469_),
    .Y(_04470_));
 sky130_fd_sc_hd__inv_1 _14871_ (.A(_12948_),
    .Y(_04471_));
 sky130_fd_sc_hd__nor3_4 _14872_ (.A(_04406_),
    .B(_12943_),
    .C(_04409_),
    .Y(_04472_));
 sky130_fd_sc_hd__o21bai_1 _14873_ (.A1(_04471_),
    .A2(_04472_),
    .B1_N(_12947_),
    .Y(_04473_));
 sky130_fd_sc_hd__a21o_4 _14874_ (.A1(_12946_),
    .A2(_04473_),
    .B1(_12945_),
    .X(_04474_));
 sky130_fd_sc_hd__xnor2_4 _14875_ (.A(_04474_),
    .B(_12952_),
    .Y(_04475_));
 sky130_fd_sc_hd__xnor2_1 _14876_ (.A(_04470_),
    .B(_04475_),
    .Y(_04476_));
 sky130_fd_sc_hd__xnor2_1 _14877_ (.A(_04467_),
    .B(_04476_),
    .Y(_12088_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1412 ();
 sky130_fd_sc_hd__or2_0 _14879_ (.A(net340),
    .B(_13241_),
    .X(\hash.CA1.S0.X[1] ));
 sky130_fd_sc_hd__inv_1 _14880_ (.A(\hash.CA1.S0.X[1] ),
    .Y(_13543_));
 sky130_fd_sc_hd__a21o_1 _14881_ (.A1(\hash.CA2.a_dash[2] ),
    .A2(_04421_),
    .B1(\hash.CA2.b_dash[2] ),
    .X(_04478_));
 sky130_fd_sc_hd__o21ai_0 _14882_ (.A1(\hash.CA2.a_dash[2] ),
    .A2(_04421_),
    .B1(_04478_),
    .Y(_12098_));
 sky130_fd_sc_hd__xnor2_2 _14883_ (.A(net1088),
    .B(net1125),
    .Y(_13246_));
 sky130_fd_sc_hd__inv_6 _14884_ (.A(_13246_),
    .Y(_12097_));
 sky130_fd_sc_hd__o21a_1 _14885_ (.A1(_12965_),
    .A2(_04419_),
    .B1(_12970_),
    .X(_04479_));
 sky130_fd_sc_hd__nor2_4 _14886_ (.A(_04479_),
    .B(_12969_),
    .Y(_04480_));
 sky130_fd_sc_hd__xor2_4 _14887_ (.A(_12968_),
    .B(_04480_),
    .X(_04481_));
 sky130_fd_sc_hd__o21a_4 _14888_ (.A1(_04433_),
    .A2(_04458_),
    .B1(_04460_),
    .X(_04482_));
 sky130_fd_sc_hd__nor2_4 _14889_ (.A(_04453_),
    .B(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__xnor2_4 _14890_ (.A(_12950_),
    .B(_04483_),
    .Y(_04484_));
 sky130_fd_sc_hd__a21o_1 _14891_ (.A1(_12924_),
    .A2(_12081_),
    .B1(_12923_),
    .X(_04485_));
 sky130_fd_sc_hd__a21oi_2 _14892_ (.A1(_12936_),
    .A2(_04485_),
    .B1(_12935_),
    .Y(_04486_));
 sky130_fd_sc_hd__xnor2_4 _14893_ (.A(_12934_),
    .B(_04486_),
    .Y(_04487_));
 sky130_fd_sc_hd__xnor2_1 _14894_ (.A(_04484_),
    .B(_04487_),
    .Y(_04488_));
 sky130_fd_sc_hd__xnor2_4 _14895_ (.A(_04488_),
    .B(_04481_),
    .Y(_12096_));
 sky130_fd_sc_hd__maj3_1 _14896_ (.A(\hash.CA2.b_dash[3] ),
    .B(\hash.CA2.a_dash[3] ),
    .C(_04470_),
    .X(_04489_));
 sky130_fd_sc_hd__inv_1 _14897_ (.A(_04489_),
    .Y(_12112_));
 sky130_fd_sc_hd__a21o_1 _14898_ (.A1(_13231_),
    .A2(_13239_),
    .B1(_13238_),
    .X(_04490_));
 sky130_fd_sc_hd__a21oi_2 _14899_ (.A1(net1125),
    .A2(_04490_),
    .B1(_13244_),
    .Y(_04491_));
 sky130_fd_sc_hd__xnor2_2 _14900_ (.A(_13252_),
    .B(_04491_),
    .Y(_13253_));
 sky130_fd_sc_hd__inv_6 _14901_ (.A(_13253_),
    .Y(_12111_));
 sky130_fd_sc_hd__clkinv_2 _14902_ (.A(_12972_),
    .Y(_04492_));
 sky130_fd_sc_hd__o21ai_2 _14903_ (.A1(_12966_),
    .A2(_12965_),
    .B1(_12970_),
    .Y(_04493_));
 sky130_fd_sc_hd__nor2_2 _14904_ (.A(_12967_),
    .B(_12969_),
    .Y(_04494_));
 sky130_fd_sc_hd__nor2_2 _14905_ (.A(_12968_),
    .B(_12967_),
    .Y(_04495_));
 sky130_fd_sc_hd__a21oi_4 _14906_ (.A1(_04493_),
    .A2(_04494_),
    .B1(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__a2111o_2 _14907_ (.A1(_04463_),
    .A2(_04465_),
    .B1(_12965_),
    .C1(_12967_),
    .D1(_12969_),
    .X(_04497_));
 sky130_fd_sc_hd__nand2_4 _14908_ (.A(_04496_),
    .B(_04497_),
    .Y(_04498_));
 sky130_fd_sc_hd__xnor2_4 _14909_ (.A(_04492_),
    .B(_04498_),
    .Y(_04499_));
 sky130_fd_sc_hd__o21ai_2 _14910_ (.A1(_04423_),
    .A2(_04424_),
    .B1(_04425_),
    .Y(_04500_));
 sky130_fd_sc_hd__xor2_4 _14911_ (.A(_12932_),
    .B(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__or2_4 _14912_ (.A(_04394_),
    .B(_04411_),
    .X(_04502_));
 sky130_fd_sc_hd__xnor2_4 _14913_ (.A(_12954_),
    .B(_04502_),
    .Y(_04503_));
 sky130_fd_sc_hd__xnor2_1 _14914_ (.A(_04501_),
    .B(_04503_),
    .Y(_04504_));
 sky130_fd_sc_hd__xnor2_2 _14915_ (.A(_04499_),
    .B(_04504_),
    .Y(_12110_));
 sky130_fd_sc_hd__maj3_1 _14916_ (.A(\hash.CA2.b_dash[4] ),
    .B(\hash.CA2.a_dash[4] ),
    .C(_04487_),
    .X(_04505_));
 sky130_fd_sc_hd__inv_1 _14917_ (.A(_04505_),
    .Y(_12121_));
 sky130_fd_sc_hd__inv_1 _14918_ (.A(_13251_),
    .Y(_04506_));
 sky130_fd_sc_hd__nor2b_2 _14919_ (.A(_12086_),
    .B_N(_13245_),
    .Y(_04507_));
 sky130_fd_sc_hd__o21ai_2 _14920_ (.A1(_13244_),
    .A2(_04507_),
    .B1(_13252_),
    .Y(_04508_));
 sky130_fd_sc_hd__a21boi_2 _14921_ (.A1(_04508_),
    .A2(_04506_),
    .B1_N(_13259_),
    .Y(_04509_));
 sky130_fd_sc_hd__nand2_1 _14922_ (.A(_04506_),
    .B(_04508_),
    .Y(_04510_));
 sky130_fd_sc_hd__nor2_2 _14923_ (.A(_13259_),
    .B(_04510_),
    .Y(_04511_));
 sky130_fd_sc_hd__nor2_4 _14924_ (.A(net1052),
    .B(_04511_),
    .Y(_13260_));
 sky130_fd_sc_hd__inv_6 _14925_ (.A(_13260_),
    .Y(_12120_));
 sky130_fd_sc_hd__o2111ai_2 _14926_ (.A1(_12965_),
    .A2(_04419_),
    .B1(_12968_),
    .C1(_12970_),
    .D1(_12972_),
    .Y(_04512_));
 sky130_fd_sc_hd__a21o_1 _14927_ (.A1(_12968_),
    .A2(_12969_),
    .B1(_12967_),
    .X(_04513_));
 sky130_fd_sc_hd__nand2_1 _14928_ (.A(_12972_),
    .B(_04513_),
    .Y(_04514_));
 sky130_fd_sc_hd__nand2_1 _14929_ (.A(_04512_),
    .B(_04514_),
    .Y(_04515_));
 sky130_fd_sc_hd__nor2_2 _14930_ (.A(_12971_),
    .B(_04515_),
    .Y(_04516_));
 sky130_fd_sc_hd__xnor2_4 _14931_ (.A(_04516_),
    .B(_12976_),
    .Y(_04517_));
 sky130_fd_sc_hd__o21ai_0 _14932_ (.A1(_04389_),
    .A2(_04436_),
    .B1(_04393_),
    .Y(_04518_));
 sky130_fd_sc_hd__a21oi_2 _14933_ (.A1(_12954_),
    .A2(_04518_),
    .B1(_12953_),
    .Y(_04519_));
 sky130_fd_sc_hd__xnor2_4 _14934_ (.A(_12956_),
    .B(_04519_),
    .Y(_04520_));
 sky130_fd_sc_hd__o21ai_2 _14935_ (.A1(_04398_),
    .A2(_04399_),
    .B1(_04400_),
    .Y(_04521_));
 sky130_fd_sc_hd__xor2_4 _14936_ (.A(_12930_),
    .B(_04521_),
    .X(_04522_));
 sky130_fd_sc_hd__xor2_1 _14937_ (.A(_04520_),
    .B(_04522_),
    .X(_04523_));
 sky130_fd_sc_hd__xnor2_2 _14938_ (.A(_04517_),
    .B(_04523_),
    .Y(_12119_));
 sky130_fd_sc_hd__maj3_1 _14939_ (.A(\hash.CA2.b_dash[5] ),
    .B(\hash.CA2.a_dash[5] ),
    .C(_04501_),
    .X(_04524_));
 sky130_fd_sc_hd__inv_2 _14940_ (.A(_04524_),
    .Y(_12130_));
 sky130_fd_sc_hd__a211oi_4 _14941_ (.A1(_13231_),
    .A2(_13239_),
    .B1(_13238_),
    .C1(_13244_),
    .Y(_04525_));
 sky130_fd_sc_hd__o211ai_1 _14942_ (.A1(_13245_),
    .A2(_13244_),
    .B1(_13252_),
    .C1(_13259_),
    .Y(_04526_));
 sky130_fd_sc_hd__a21oi_2 _14943_ (.A1(_13259_),
    .A2(_13251_),
    .B1(_13258_),
    .Y(_04527_));
 sky130_fd_sc_hd__o21ai_4 _14944_ (.A1(_04525_),
    .A2(_04526_),
    .B1(_04527_),
    .Y(_04528_));
 sky130_fd_sc_hd__xor2_2 _14945_ (.A(_13266_),
    .B(_04528_),
    .X(_13267_));
 sky130_fd_sc_hd__inv_6 _14946_ (.A(_13267_),
    .Y(_12129_));
 sky130_fd_sc_hd__nor2_1 _14947_ (.A(_04492_),
    .B(_04498_),
    .Y(_04529_));
 sky130_fd_sc_hd__o21ai_1 _14948_ (.A1(_12971_),
    .A2(_04529_),
    .B1(_12976_),
    .Y(_04530_));
 sky130_fd_sc_hd__nor2_1 _14949_ (.A(_12974_),
    .B(_12975_),
    .Y(_04531_));
 sky130_fd_sc_hd__and3_4 _14950_ (.A(_12974_),
    .B(_12972_),
    .C(_12976_),
    .X(_04532_));
 sky130_fd_sc_hd__nand3_4 _14951_ (.A(_04496_),
    .B(_04497_),
    .C(_04532_),
    .Y(_04533_));
 sky130_fd_sc_hd__nand2_4 _14952_ (.A(_12974_),
    .B(_12975_),
    .Y(_04534_));
 sky130_fd_sc_hd__nand3_4 _14953_ (.A(_12974_),
    .B(_12976_),
    .C(_12971_),
    .Y(_04535_));
 sky130_fd_sc_hd__nand3_4 _14954_ (.A(_04533_),
    .B(_04534_),
    .C(_04535_),
    .Y(_04536_));
 sky130_fd_sc_hd__a21oi_4 _14955_ (.A1(_04530_),
    .A2(_04531_),
    .B1(_04536_),
    .Y(_04537_));
 sky130_fd_sc_hd__nor2_1 _14956_ (.A(_04394_),
    .B(_04411_),
    .Y(_04538_));
 sky130_fd_sc_hd__a21o_1 _14957_ (.A1(_12954_),
    .A2(_04538_),
    .B1(_12953_),
    .X(_04539_));
 sky130_fd_sc_hd__a21oi_2 _14958_ (.A1(_12956_),
    .A2(_04539_),
    .B1(_12955_),
    .Y(_04540_));
 sky130_fd_sc_hd__xnor2_4 _14959_ (.A(_12958_),
    .B(_04540_),
    .Y(_04541_));
 sky130_fd_sc_hd__xnor2_4 _14960_ (.A(_12928_),
    .B(_04428_),
    .Y(_04542_));
 sky130_fd_sc_hd__inv_6 _14961_ (.A(_04542_),
    .Y(_04543_));
 sky130_fd_sc_hd__xnor2_1 _14962_ (.A(_04541_),
    .B(_04543_),
    .Y(_04544_));
 sky130_fd_sc_hd__xnor2_2 _14963_ (.A(_04537_),
    .B(_04544_),
    .Y(_12128_));
 sky130_fd_sc_hd__maj3_1 _14964_ (.A(\hash.CA2.b_dash[6] ),
    .B(\hash.CA2.a_dash[6] ),
    .C(_04522_),
    .X(_04545_));
 sky130_fd_sc_hd__inv_2 _14965_ (.A(_04545_),
    .Y(_12139_));
 sky130_fd_sc_hd__o21a_1 _14966_ (.A1(_04509_),
    .A2(_13258_),
    .B1(_13266_),
    .X(_04546_));
 sky130_fd_sc_hd__or2_4 _14967_ (.A(_13265_),
    .B(_04546_),
    .X(_04547_));
 sky130_fd_sc_hd__xor2_4 _14968_ (.A(_13273_),
    .B(_04547_),
    .X(_13274_));
 sky130_fd_sc_hd__inv_4 _14969_ (.A(_13274_),
    .Y(_12138_));
 sky130_fd_sc_hd__nor3_1 _14970_ (.A(_12971_),
    .B(_12973_),
    .C(_12975_),
    .Y(_04548_));
 sky130_fd_sc_hd__nand3_2 _14971_ (.A(_04512_),
    .B(_04514_),
    .C(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hd__nor3_1 _14972_ (.A(_12976_),
    .B(_12973_),
    .C(_12975_),
    .Y(_04550_));
 sky130_fd_sc_hd__nor2_1 _14973_ (.A(_12974_),
    .B(_12973_),
    .Y(_04551_));
 sky130_fd_sc_hd__nor2_2 _14974_ (.A(_04550_),
    .B(_04551_),
    .Y(_04552_));
 sky130_fd_sc_hd__nand2_4 _14975_ (.A(_04549_),
    .B(_04552_),
    .Y(_04553_));
 sky130_fd_sc_hd__xnor2_4 _14976_ (.A(_04553_),
    .B(_12978_),
    .Y(_04554_));
 sky130_fd_sc_hd__nor2_1 _14977_ (.A(_04455_),
    .B(_04483_),
    .Y(_04555_));
 sky130_fd_sc_hd__a22o_1 _14978_ (.A1(_12964_),
    .A2(_04450_),
    .B1(_04453_),
    .B2(_04456_),
    .X(_04556_));
 sky130_fd_sc_hd__and2_4 _14979_ (.A(_04482_),
    .B(_04456_),
    .X(_04557_));
 sky130_fd_sc_hd__nor2_1 _14980_ (.A(_04556_),
    .B(_04557_),
    .Y(_04558_));
 sky130_fd_sc_hd__o31a_1 _14981_ (.A1(_12964_),
    .A2(_04450_),
    .A3(_04555_),
    .B1(_04558_),
    .X(_04559_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1411 ();
 sky130_fd_sc_hd__nand2_2 _14983_ (.A(_04397_),
    .B(net1085),
    .Y(_04561_));
 sky130_fd_sc_hd__xnor2_4 _14984_ (.A(_12940_),
    .B(_04561_),
    .Y(_04562_));
 sky130_fd_sc_hd__xor2_1 _14985_ (.A(_04559_),
    .B(_04562_),
    .X(_04563_));
 sky130_fd_sc_hd__xnor2_2 _14986_ (.A(_04554_),
    .B(_04563_),
    .Y(_12137_));
 sky130_fd_sc_hd__maj3_1 _14987_ (.A(\hash.CA2.b_dash[7] ),
    .B(\hash.CA2.a_dash[7] ),
    .C(_04542_),
    .X(_04564_));
 sky130_fd_sc_hd__inv_1 _14988_ (.A(_04564_),
    .Y(_12148_));
 sky130_fd_sc_hd__clkinv_1 _14989_ (.A(_13272_),
    .Y(_04565_));
 sky130_fd_sc_hd__o21ai_0 _14990_ (.A1(_13266_),
    .A2(_13265_),
    .B1(_13273_),
    .Y(_04566_));
 sky130_fd_sc_hd__nand2_1 _14991_ (.A(_04565_),
    .B(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__o31ai_2 _14992_ (.A1(_13265_),
    .A2(_13272_),
    .A3(_04528_),
    .B1(_04567_),
    .Y(_04568_));
 sky130_fd_sc_hd__xnor2_2 _14993_ (.A(_13280_),
    .B(_04568_),
    .Y(_13281_));
 sky130_fd_sc_hd__inv_4 _14994_ (.A(_13281_),
    .Y(_12147_));
 sky130_fd_sc_hd__o21ai_2 _14995_ (.A1(_12973_),
    .A2(_04536_),
    .B1(_12978_),
    .Y(_04569_));
 sky130_fd_sc_hd__nor2_2 _14996_ (.A(_12980_),
    .B(_12977_),
    .Y(_04570_));
 sky130_fd_sc_hd__nor2_2 _14997_ (.A(_12973_),
    .B(_12977_),
    .Y(_04571_));
 sky130_fd_sc_hd__o21ai_2 _14998_ (.A1(_12978_),
    .A2(_12977_),
    .B1(_12980_),
    .Y(_04572_));
 sky130_fd_sc_hd__a41oi_4 _14999_ (.A1(_04533_),
    .A2(_04534_),
    .A3(_04535_),
    .A4(_04571_),
    .B1(_04572_),
    .Y(_04573_));
 sky130_fd_sc_hd__a21o_4 _15000_ (.A1(_04569_),
    .A2(_04570_),
    .B1(_04573_),
    .X(_04574_));
 sky130_fd_sc_hd__o21ai_0 _15001_ (.A1(_04502_),
    .A2(_04412_),
    .B1(_04383_),
    .Y(_04575_));
 sky130_fd_sc_hd__a21o_4 _15002_ (.A1(_12964_),
    .A2(_04575_),
    .B1(_12963_),
    .X(_04576_));
 sky130_fd_sc_hd__xor2_2 _15003_ (.A(_12962_),
    .B(_04576_),
    .X(_04577_));
 sky130_fd_sc_hd__a21o_1 _15004_ (.A1(_12940_),
    .A2(_12927_),
    .B1(_12939_),
    .X(_04578_));
 sky130_fd_sc_hd__a41oi_2 _15005_ (.A1(_12928_),
    .A2(_12940_),
    .A3(_04422_),
    .A4(_04427_),
    .B1(_04578_),
    .Y(_04579_));
 sky130_fd_sc_hd__xnor2_4 _15006_ (.A(_12938_),
    .B(_04579_),
    .Y(_04580_));
 sky130_fd_sc_hd__xnor2_1 _15007_ (.A(_04577_),
    .B(_04580_),
    .Y(_04581_));
 sky130_fd_sc_hd__xnor2_2 _15008_ (.A(_04574_),
    .B(_04581_),
    .Y(_12146_));
 sky130_fd_sc_hd__maj3_1 _15009_ (.A(\hash.CA2.b_dash[8] ),
    .B(\hash.CA2.a_dash[8] ),
    .C(_04562_),
    .X(_04582_));
 sky130_fd_sc_hd__inv_2 _15010_ (.A(_04582_),
    .Y(_12157_));
 sky130_fd_sc_hd__o21ai_2 _15011_ (.A1(_13265_),
    .A2(_04546_),
    .B1(_13273_),
    .Y(_04583_));
 sky130_fd_sc_hd__nand2_1 _15012_ (.A(_04565_),
    .B(_04583_),
    .Y(_04584_));
 sky130_fd_sc_hd__a21o_1 _15013_ (.A1(_04584_),
    .A2(_13280_),
    .B1(_13279_),
    .X(_04585_));
 sky130_fd_sc_hd__xor2_4 _15014_ (.A(_13287_),
    .B(_04585_),
    .X(_13288_));
 sky130_fd_sc_hd__inv_4 _15015_ (.A(_13288_),
    .Y(_12156_));
 sky130_fd_sc_hd__a31o_1 _15016_ (.A1(_12978_),
    .A2(_04549_),
    .A3(_04552_),
    .B1(_12977_),
    .X(_04586_));
 sky130_fd_sc_hd__a21oi_4 _15017_ (.A1(_12980_),
    .A2(_04586_),
    .B1(_12979_),
    .Y(_04587_));
 sky130_fd_sc_hd__xor2_4 _15018_ (.A(_12982_),
    .B(_04587_),
    .X(_04588_));
 sky130_fd_sc_hd__clkinv_1 _15019_ (.A(_12960_),
    .Y(_04589_));
 sky130_fd_sc_hd__nor3_1 _15020_ (.A(_04589_),
    .B(_12961_),
    .C(_12963_),
    .Y(_04590_));
 sky130_fd_sc_hd__nand2_2 _15021_ (.A(_04558_),
    .B(_04590_),
    .Y(_04591_));
 sky130_fd_sc_hd__nor2b_4 _15022_ (.A(_12960_),
    .B_N(_12962_),
    .Y(_04592_));
 sky130_fd_sc_hd__o21ai_2 _15023_ (.A1(_04556_),
    .A2(_04557_),
    .B1(_04592_),
    .Y(_04593_));
 sky130_fd_sc_hd__nor3_1 _15024_ (.A(_04589_),
    .B(_12962_),
    .C(_12961_),
    .Y(_04594_));
 sky130_fd_sc_hd__a221oi_2 _15025_ (.A1(_04589_),
    .A2(_12961_),
    .B1(_12963_),
    .B2(_04592_),
    .C1(_04594_),
    .Y(_04595_));
 sky130_fd_sc_hd__nand3_4 _15026_ (.A(_04591_),
    .B(_04593_),
    .C(_04595_),
    .Y(_04596_));
 sky130_fd_sc_hd__a31o_1 _15027_ (.A1(_12940_),
    .A2(_04397_),
    .A3(_04402_),
    .B1(_12939_),
    .X(_04597_));
 sky130_fd_sc_hd__a21oi_2 _15028_ (.A1(_12938_),
    .A2(_04597_),
    .B1(_12937_),
    .Y(_04598_));
 sky130_fd_sc_hd__xnor2_4 _15029_ (.A(_12942_),
    .B(_04598_),
    .Y(_04599_));
 sky130_fd_sc_hd__xnor2_1 _15030_ (.A(_04596_),
    .B(_04599_),
    .Y(_04600_));
 sky130_fd_sc_hd__xnor2_4 _15031_ (.A(_04600_),
    .B(net1095),
    .Y(_12155_));
 sky130_fd_sc_hd__maj3_1 _15032_ (.A(\hash.CA2.b_dash[9] ),
    .B(\hash.CA2.a_dash[9] ),
    .C(_04580_),
    .X(_04601_));
 sky130_fd_sc_hd__inv_4 _15033_ (.A(_04601_),
    .Y(_12166_));
 sky130_fd_sc_hd__nor2b_1 _15034_ (.A(_04568_),
    .B_N(_13280_),
    .Y(_04602_));
 sky130_fd_sc_hd__o21ai_0 _15035_ (.A1(_13279_),
    .A2(_04602_),
    .B1(_13287_),
    .Y(_04603_));
 sky130_fd_sc_hd__nand2b_2 _15036_ (.A_N(_13286_),
    .B(_04603_),
    .Y(_04604_));
 sky130_fd_sc_hd__xor2_2 _15037_ (.A(_13294_),
    .B(_04604_),
    .X(_13295_));
 sky130_fd_sc_hd__inv_4 _15038_ (.A(_13295_),
    .Y(_12165_));
 sky130_fd_sc_hd__xor2_1 _15039_ (.A(\hash.CA2.p1[31] ),
    .B(\hash.CA2.p3[31] ),
    .X(_04605_));
 sky130_fd_sc_hd__or3_1 _15040_ (.A(_12979_),
    .B(_12981_),
    .C(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__nand2_1 _15041_ (.A(_12982_),
    .B(_04605_),
    .Y(_04607_));
 sky130_fd_sc_hd__mux2i_2 _15042_ (.A0(_04606_),
    .A1(_04607_),
    .S(_04573_),
    .Y(_04608_));
 sky130_fd_sc_hd__and2_0 _15043_ (.A(_12982_),
    .B(_12979_),
    .X(_04609_));
 sky130_fd_sc_hd__o21ai_0 _15044_ (.A1(_12981_),
    .A2(_04609_),
    .B1(_04605_),
    .Y(_04610_));
 sky130_fd_sc_hd__o31ai_2 _15045_ (.A1(_12982_),
    .A2(_12981_),
    .A3(_04605_),
    .B1(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__nor2_4 _15046_ (.A(_04611_),
    .B(_04608_),
    .Y(_04612_));
 sky130_fd_sc_hd__nor2_2 _15047_ (.A(_04433_),
    .B(_04458_),
    .Y(_04613_));
 sky130_fd_sc_hd__xnor2_4 _15048_ (.A(_12944_),
    .B(_04613_),
    .Y(_04614_));
 sky130_fd_sc_hd__xor2_1 _15049_ (.A(_04420_),
    .B(_04614_),
    .X(_04615_));
 sky130_fd_sc_hd__xnor2_2 _15050_ (.A(_04612_),
    .B(_04615_),
    .Y(_12164_));
 sky130_fd_sc_hd__maj3_1 _15051_ (.A(\hash.CA2.b_dash[10] ),
    .B(\hash.CA2.a_dash[10] ),
    .C(_04599_),
    .X(_04616_));
 sky130_fd_sc_hd__clkinv_2 _15052_ (.A(_04616_),
    .Y(_12175_));
 sky130_fd_sc_hd__and3_1 _15053_ (.A(_13280_),
    .B(_13287_),
    .C(_13294_),
    .X(_04617_));
 sky130_fd_sc_hd__a21boi_2 _15054_ (.A1(_04583_),
    .A2(_04565_),
    .B1_N(_04617_),
    .Y(_04618_));
 sky130_fd_sc_hd__a21oi_4 _15055_ (.A1(_13287_),
    .A2(_13279_),
    .B1(_13286_),
    .Y(_04619_));
 sky130_fd_sc_hd__nor2b_4 _15056_ (.A(_04619_),
    .B_N(_13294_),
    .Y(_04620_));
 sky130_fd_sc_hd__nor2_1 _15057_ (.A(_13293_),
    .B(_04620_),
    .Y(_04621_));
 sky130_fd_sc_hd__nand2b_1 _15058_ (.A_N(_04618_),
    .B(_04621_),
    .Y(_04622_));
 sky130_fd_sc_hd__xor2_1 _15059_ (.A(_13301_),
    .B(_04622_),
    .X(_13302_));
 sky130_fd_sc_hd__inv_4 _15060_ (.A(_13302_),
    .Y(_12174_));
 sky130_fd_sc_hd__xnor2_4 _15061_ (.A(_12948_),
    .B(_04472_),
    .Y(_04623_));
 sky130_fd_sc_hd__xnor2_1 _15062_ (.A(_12922_),
    .B(_04623_),
    .Y(_04624_));
 sky130_fd_sc_hd__xor2_1 _15063_ (.A(_04467_),
    .B(_04624_),
    .X(_12173_));
 sky130_fd_sc_hd__maj3_1 _15064_ (.A(\hash.CA2.b_dash[11] ),
    .B(\hash.CA2.a_dash[11] ),
    .C(_04614_),
    .X(_04625_));
 sky130_fd_sc_hd__inv_1 _15065_ (.A(_04625_),
    .Y(_12184_));
 sky130_fd_sc_hd__o311ai_4 _15066_ (.A1(_13265_),
    .A2(_13272_),
    .A3(_04528_),
    .B1(_04567_),
    .C1(_04617_),
    .Y(_04626_));
 sky130_fd_sc_hd__a21boi_2 _15067_ (.A1(_04626_),
    .A2(_04621_),
    .B1_N(_13301_),
    .Y(_04627_));
 sky130_fd_sc_hd__nor2_1 _15068_ (.A(_13300_),
    .B(_04627_),
    .Y(_04628_));
 sky130_fd_sc_hd__xnor2_2 _15069_ (.A(_13308_),
    .B(_04628_),
    .Y(_13309_));
 sky130_fd_sc_hd__inv_4 _15070_ (.A(_13309_),
    .Y(_12183_));
 sky130_fd_sc_hd__xnor2_1 _15071_ (.A(_12082_),
    .B(_04437_),
    .Y(_04629_));
 sky130_fd_sc_hd__xnor2_1 _15072_ (.A(_04481_),
    .B(_04629_),
    .Y(_12182_));
 sky130_fd_sc_hd__maj3_4 _15073_ (.A(\hash.CA2.b_dash[12] ),
    .B(\hash.CA2.a_dash[12] ),
    .C(_04623_),
    .X(_04630_));
 sky130_fd_sc_hd__inv_1 _15074_ (.A(_04630_),
    .Y(_12193_));
 sky130_fd_sc_hd__or3_4 _15075_ (.A(_13293_),
    .B(_13300_),
    .C(_13307_),
    .X(_04631_));
 sky130_fd_sc_hd__nor3_1 _15076_ (.A(_13301_),
    .B(_13300_),
    .C(_13307_),
    .Y(_04632_));
 sky130_fd_sc_hd__nor2_1 _15077_ (.A(_13308_),
    .B(_13307_),
    .Y(_04633_));
 sky130_fd_sc_hd__nor2_2 _15078_ (.A(_04632_),
    .B(_04633_),
    .Y(_04634_));
 sky130_fd_sc_hd__o31ai_4 _15079_ (.A1(_04620_),
    .A2(_04631_),
    .A3(_04618_),
    .B1(_04634_),
    .Y(_04635_));
 sky130_fd_sc_hd__xnor2_4 _15080_ (.A(_13315_),
    .B(net1053),
    .Y(_13316_));
 sky130_fd_sc_hd__inv_4 _15081_ (.A(_13316_),
    .Y(_12192_));
 sky130_fd_sc_hd__xor2_2 _15082_ (.A(_12952_),
    .B(_04474_),
    .X(_04636_));
 sky130_fd_sc_hd__xnor2_1 _15083_ (.A(_04421_),
    .B(_04636_),
    .Y(_04637_));
 sky130_fd_sc_hd__xnor2_1 _15084_ (.A(_04499_),
    .B(_04637_),
    .Y(_12191_));
 sky130_fd_sc_hd__nor2_2 _15085_ (.A(\hash.CA2.a_dash[13] ),
    .B(_04437_),
    .Y(_04638_));
 sky130_fd_sc_hd__a21oi_1 _15086_ (.A1(\hash.CA2.a_dash[13] ),
    .A2(_04437_),
    .B1(\hash.CA2.b_dash[13] ),
    .Y(_04639_));
 sky130_fd_sc_hd__nor2_1 _15087_ (.A(_04638_),
    .B(_04639_),
    .Y(_04640_));
 sky130_fd_sc_hd__clkinv_1 _15088_ (.A(_04640_),
    .Y(_12202_));
 sky130_fd_sc_hd__clkinv_2 _15089_ (.A(_13322_),
    .Y(_04641_));
 sky130_fd_sc_hd__o21ai_1 _15090_ (.A1(_04627_),
    .A2(_13300_),
    .B1(_13308_),
    .Y(_04642_));
 sky130_fd_sc_hd__nand2b_1 _15091_ (.A_N(_13307_),
    .B(_04642_),
    .Y(_04643_));
 sky130_fd_sc_hd__a21o_1 _15092_ (.A1(_04643_),
    .A2(_13315_),
    .B1(_13314_),
    .X(_04644_));
 sky130_fd_sc_hd__xnor2_2 _15093_ (.A(_04641_),
    .B(_04644_),
    .Y(_13323_));
 sky130_fd_sc_hd__inv_4 _15094_ (.A(_13323_),
    .Y(_12201_));
 sky130_fd_sc_hd__xor2_1 _15095_ (.A(_04470_),
    .B(_04484_),
    .X(_04645_));
 sky130_fd_sc_hd__xnor2_1 _15096_ (.A(_04517_),
    .B(_04645_),
    .Y(_12200_));
 sky130_fd_sc_hd__nor2_1 _15097_ (.A(\hash.CA2.a_dash[14] ),
    .B(_04636_),
    .Y(_04646_));
 sky130_fd_sc_hd__a21oi_1 _15098_ (.A1(\hash.CA2.a_dash[14] ),
    .A2(_04636_),
    .B1(\hash.CA2.b_dash[14] ),
    .Y(_04647_));
 sky130_fd_sc_hd__nor2_1 _15099_ (.A(_04646_),
    .B(_04647_),
    .Y(_04648_));
 sky130_fd_sc_hd__inv_1 _15100_ (.A(_04648_),
    .Y(_12211_));
 sky130_fd_sc_hd__inv_1 _15101_ (.A(_13315_),
    .Y(_04649_));
 sky130_fd_sc_hd__nor2_1 _15102_ (.A(_04649_),
    .B(_04641_),
    .Y(_04650_));
 sky130_fd_sc_hd__nand2_1 _15103_ (.A(_13329_),
    .B(_04650_),
    .Y(_04651_));
 sky130_fd_sc_hd__and3_1 _15104_ (.A(_13322_),
    .B(_13329_),
    .C(_13314_),
    .X(_04652_));
 sky130_fd_sc_hd__a21oi_2 _15105_ (.A1(_13329_),
    .A2(_13321_),
    .B1(_04652_),
    .Y(_04653_));
 sky130_fd_sc_hd__o21ai_4 _15106_ (.A1(net1053),
    .A2(_04651_),
    .B1(_04653_),
    .Y(_04654_));
 sky130_fd_sc_hd__o21bai_1 _15107_ (.A1(_04649_),
    .A2(_04635_),
    .B1_N(_13314_),
    .Y(_04655_));
 sky130_fd_sc_hd__a211oi_1 _15108_ (.A1(_13322_),
    .A2(_04655_),
    .B1(_13321_),
    .C1(_13329_),
    .Y(_04656_));
 sky130_fd_sc_hd__nor2_2 _15109_ (.A(_04656_),
    .B(_04654_),
    .Y(_13330_));
 sky130_fd_sc_hd__inv_4 _15110_ (.A(net1050),
    .Y(_12210_));
 sky130_fd_sc_hd__xor2_1 _15111_ (.A(_04487_),
    .B(_04503_),
    .X(_04657_));
 sky130_fd_sc_hd__xnor2_1 _15112_ (.A(net1072),
    .B(_04657_),
    .Y(_12209_));
 sky130_fd_sc_hd__maj3_1 _15113_ (.A(\hash.CA2.b_dash[15] ),
    .B(\hash.CA2.a_dash[15] ),
    .C(_04484_),
    .X(_04658_));
 sky130_fd_sc_hd__inv_1 _15114_ (.A(_04658_),
    .Y(_12220_));
 sky130_fd_sc_hd__a211oi_2 _15115_ (.A1(_04644_),
    .A2(_13322_),
    .B1(_13328_),
    .C1(_13321_),
    .Y(_04659_));
 sky130_fd_sc_hd__nor2_1 _15116_ (.A(_13329_),
    .B(_13328_),
    .Y(_04660_));
 sky130_fd_sc_hd__nor2_4 _15117_ (.A(_04660_),
    .B(_04659_),
    .Y(_04661_));
 sky130_fd_sc_hd__xor2_2 _15118_ (.A(_13336_),
    .B(_04661_),
    .X(_13337_));
 sky130_fd_sc_hd__inv_4 _15119_ (.A(_13337_),
    .Y(_12219_));
 sky130_fd_sc_hd__xor2_4 _15120_ (.A(_12978_),
    .B(_04553_),
    .X(_04662_));
 sky130_fd_sc_hd__xnor2_1 _15121_ (.A(_04501_),
    .B(_04520_),
    .Y(_04663_));
 sky130_fd_sc_hd__xnor2_1 _15122_ (.A(_04662_),
    .B(_04663_),
    .Y(_12218_));
 sky130_fd_sc_hd__maj3_1 _15123_ (.A(\hash.CA2.b_dash[16] ),
    .B(\hash.CA2.a_dash[16] ),
    .C(_04503_),
    .X(_04664_));
 sky130_fd_sc_hd__clkinvlp_2 _15124_ (.A(_04664_),
    .Y(_12229_));
 sky130_fd_sc_hd__o21ai_1 _15125_ (.A1(_13328_),
    .A2(_04654_),
    .B1(_13336_),
    .Y(_04665_));
 sky130_fd_sc_hd__nand2b_2 _15126_ (.A_N(_13335_),
    .B(_04665_),
    .Y(_04666_));
 sky130_fd_sc_hd__xor2_4 _15127_ (.A(_13343_),
    .B(_04666_),
    .X(_13344_));
 sky130_fd_sc_hd__inv_4 _15128_ (.A(net1099),
    .Y(_12228_));
 sky130_fd_sc_hd__xnor2_1 _15129_ (.A(_04522_),
    .B(_04541_),
    .Y(_04667_));
 sky130_fd_sc_hd__xnor2_1 _15130_ (.A(_04574_),
    .B(_04667_),
    .Y(_12227_));
 sky130_fd_sc_hd__maj3_1 _15131_ (.A(\hash.CA2.b_dash[17] ),
    .B(\hash.CA2.a_dash[17] ),
    .C(_04520_),
    .X(_04668_));
 sky130_fd_sc_hd__inv_2 _15132_ (.A(_04668_),
    .Y(_12238_));
 sky130_fd_sc_hd__a21o_1 _15133_ (.A1(_13336_),
    .A2(_04661_),
    .B1(_13335_),
    .X(_04669_));
 sky130_fd_sc_hd__a21o_1 _15134_ (.A1(_13343_),
    .A2(_04669_),
    .B1(_13342_),
    .X(_04670_));
 sky130_fd_sc_hd__xor2_2 _15135_ (.A(_13350_),
    .B(_04670_),
    .X(_13351_));
 sky130_fd_sc_hd__inv_4 _15136_ (.A(net1065),
    .Y(_12237_));
 sky130_fd_sc_hd__xnor2_1 _15137_ (.A(_04542_),
    .B(_04559_),
    .Y(_04671_));
 sky130_fd_sc_hd__xnor2_2 _15138_ (.A(net1095),
    .B(_04671_),
    .Y(_12236_));
 sky130_fd_sc_hd__nor2_1 _15139_ (.A(\hash.CA2.a_dash[18] ),
    .B(_04541_),
    .Y(_04672_));
 sky130_fd_sc_hd__a21oi_1 _15140_ (.A1(\hash.CA2.a_dash[18] ),
    .A2(_04541_),
    .B1(\hash.CA2.b_dash[18] ),
    .Y(_04673_));
 sky130_fd_sc_hd__nor2_2 _15141_ (.A(_04672_),
    .B(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__inv_1 _15142_ (.A(_04674_),
    .Y(_12247_));
 sky130_fd_sc_hd__a21o_1 _15143_ (.A1(_13336_),
    .A2(_13328_),
    .B1(_13335_),
    .X(_04675_));
 sky130_fd_sc_hd__a21o_1 _15144_ (.A1(_13343_),
    .A2(_04675_),
    .B1(_13342_),
    .X(_04676_));
 sky130_fd_sc_hd__a21oi_1 _15145_ (.A1(_13350_),
    .A2(_04676_),
    .B1(_13349_),
    .Y(_04677_));
 sky130_fd_sc_hd__and3_4 _15146_ (.A(_13336_),
    .B(_13343_),
    .C(_13350_),
    .X(_04678_));
 sky130_fd_sc_hd__nand2_1 _15147_ (.A(_04654_),
    .B(_04678_),
    .Y(_04679_));
 sky130_fd_sc_hd__nand2_1 _15148_ (.A(_04677_),
    .B(_04679_),
    .Y(_04680_));
 sky130_fd_sc_hd__xor2_2 _15149_ (.A(_13357_),
    .B(_04680_),
    .X(_13358_));
 sky130_fd_sc_hd__inv_4 _15150_ (.A(_13358_),
    .Y(_12246_));
 sky130_fd_sc_hd__xnor2_2 _15151_ (.A(_12962_),
    .B(_04576_),
    .Y(_04681_));
 sky130_fd_sc_hd__xnor2_1 _15152_ (.A(_04562_),
    .B(_04681_),
    .Y(_04682_));
 sky130_fd_sc_hd__xnor2_1 _15153_ (.A(_04612_),
    .B(_04682_),
    .Y(_12245_));
 sky130_fd_sc_hd__maj3_4 _15154_ (.A(\hash.CA2.b_dash[19] ),
    .B(\hash.CA2.a_dash[19] ),
    .C(_04559_),
    .X(_04683_));
 sky130_fd_sc_hd__inv_1 _15155_ (.A(_04683_),
    .Y(_12256_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1410 ();
 sky130_fd_sc_hd__a21o_1 _15157_ (.A1(_13343_),
    .A2(_13335_),
    .B1(_13342_),
    .X(_04685_));
 sky130_fd_sc_hd__a21o_1 _15158_ (.A1(_13350_),
    .A2(_04685_),
    .B1(_13349_),
    .X(_04686_));
 sky130_fd_sc_hd__a21o_4 _15159_ (.A1(_13357_),
    .A2(_04686_),
    .B1(_13356_),
    .X(_04687_));
 sky130_fd_sc_hd__a31oi_4 _15160_ (.A1(_13357_),
    .A2(_04661_),
    .A3(_04678_),
    .B1(_04687_),
    .Y(_04688_));
 sky130_fd_sc_hd__xnor2_2 _15161_ (.A(_13364_),
    .B(net1090),
    .Y(_13365_));
 sky130_fd_sc_hd__inv_4 _15162_ (.A(_13365_),
    .Y(_12255_));
 sky130_fd_sc_hd__xnor2_1 _15163_ (.A(_12922_),
    .B(_04580_),
    .Y(_04689_));
 sky130_fd_sc_hd__xor2_1 _15164_ (.A(_04596_),
    .B(_04689_),
    .X(_12254_));
 sky130_fd_sc_hd__maj3_1 _15165_ (.A(\hash.CA2.b_dash[20] ),
    .B(\hash.CA2.a_dash[20] ),
    .C(_04577_),
    .X(_04690_));
 sky130_fd_sc_hd__clkinv_2 _15166_ (.A(_04690_),
    .Y(_12265_));
 sky130_fd_sc_hd__nand2_1 _15167_ (.A(_13357_),
    .B(_13364_),
    .Y(_04691_));
 sky130_fd_sc_hd__nand2_1 _15168_ (.A(_13364_),
    .B(_13356_),
    .Y(_04692_));
 sky130_fd_sc_hd__o21ai_0 _15169_ (.A1(_04677_),
    .A2(_04691_),
    .B1(_04692_),
    .Y(_04693_));
 sky130_fd_sc_hd__a41oi_2 _15170_ (.A1(_13357_),
    .A2(_13364_),
    .A3(_04654_),
    .A4(_04678_),
    .B1(_04693_),
    .Y(_04694_));
 sky130_fd_sc_hd__nor2b_1 _15171_ (.A(_13363_),
    .B_N(_04694_),
    .Y(_04695_));
 sky130_fd_sc_hd__xnor2_2 _15172_ (.A(_13371_),
    .B(_04695_),
    .Y(_13372_));
 sky130_fd_sc_hd__inv_4 _15173_ (.A(_13372_),
    .Y(_12264_));
 sky130_fd_sc_hd__xnor2_1 _15174_ (.A(_12082_),
    .B(_04599_),
    .Y(_04696_));
 sky130_fd_sc_hd__xor2_1 _15175_ (.A(_04420_),
    .B(_04696_),
    .X(_12263_));
 sky130_fd_sc_hd__nor2_2 _15176_ (.A(\hash.CA2.a_dash[21] ),
    .B(_04596_),
    .Y(_04697_));
 sky130_fd_sc_hd__a21oi_1 _15177_ (.A1(\hash.CA2.a_dash[21] ),
    .A2(_04596_),
    .B1(\hash.CA2.b_dash[21] ),
    .Y(_04698_));
 sky130_fd_sc_hd__nor2_1 _15178_ (.A(_04697_),
    .B(_04698_),
    .Y(_04699_));
 sky130_fd_sc_hd__clkinv_1 _15179_ (.A(_04699_),
    .Y(_12274_));
 sky130_fd_sc_hd__inv_1 _15180_ (.A(_13364_),
    .Y(_04700_));
 sky130_fd_sc_hd__o21bai_1 _15181_ (.A1(_04688_),
    .A2(_04700_),
    .B1_N(_13363_),
    .Y(_04701_));
 sky130_fd_sc_hd__a21oi_2 _15182_ (.A1(_13371_),
    .A2(_04701_),
    .B1(_13370_),
    .Y(_04702_));
 sky130_fd_sc_hd__xnor2_2 _15183_ (.A(_13378_),
    .B(_04702_),
    .Y(_13379_));
 sky130_fd_sc_hd__clkinvlp_2 _15184_ (.A(net1068),
    .Y(_12273_));
 sky130_fd_sc_hd__xor2_1 _15185_ (.A(_04421_),
    .B(_04614_),
    .X(_04703_));
 sky130_fd_sc_hd__xnor2_1 _15186_ (.A(_04467_),
    .B(_04703_),
    .Y(_12272_));
 sky130_fd_sc_hd__nand2_2 _15187_ (.A(\hash.CA2.a_dash[22] ),
    .B(_04420_),
    .Y(_04704_));
 sky130_fd_sc_hd__o21ai_0 _15188_ (.A1(\hash.CA2.a_dash[22] ),
    .A2(_04420_),
    .B1(\hash.CA2.b_dash[22] ),
    .Y(_04705_));
 sky130_fd_sc_hd__nand2_2 _15189_ (.A(_04704_),
    .B(_04705_),
    .Y(_04706_));
 sky130_fd_sc_hd__inv_2 _15190_ (.A(_04706_),
    .Y(_12283_));
 sky130_fd_sc_hd__nor3_2 _15191_ (.A(_13363_),
    .B(_13370_),
    .C(_13377_),
    .Y(_04707_));
 sky130_fd_sc_hd__or2_4 _15192_ (.A(_13371_),
    .B(_13370_),
    .X(_04708_));
 sky130_fd_sc_hd__a21oi_2 _15193_ (.A1(_13378_),
    .A2(_04708_),
    .B1(_13377_),
    .Y(_04709_));
 sky130_fd_sc_hd__a21oi_4 _15194_ (.A1(_04694_),
    .A2(_04707_),
    .B1(_04709_),
    .Y(_04710_));
 sky130_fd_sc_hd__xor2_4 _15195_ (.A(_13385_),
    .B(net1051),
    .X(_13386_));
 sky130_fd_sc_hd__clkinvlp_2 _15196_ (.A(net1067),
    .Y(_12282_));
 sky130_fd_sc_hd__xnor2_1 _15197_ (.A(_04470_),
    .B(_04623_),
    .Y(_04711_));
 sky130_fd_sc_hd__xnor2_2 _15198_ (.A(net1107),
    .B(_04711_),
    .Y(_12281_));
 sky130_fd_sc_hd__maj3_1 _15199_ (.A(\hash.CA2.b_dash[23] ),
    .B(\hash.CA2.a_dash[23] ),
    .C(_04467_),
    .X(_04712_));
 sky130_fd_sc_hd__inv_4 _15200_ (.A(_04712_),
    .Y(_12292_));
 sky130_fd_sc_hd__a211o_1 _15201_ (.A1(_13364_),
    .A2(_04687_),
    .B1(_13370_),
    .C1(_13363_),
    .X(_04713_));
 sky130_fd_sc_hd__and3_1 _15202_ (.A(_13378_),
    .B(_13385_),
    .C(_04708_),
    .X(_04714_));
 sky130_fd_sc_hd__a221oi_1 _15203_ (.A1(_13385_),
    .A2(_13377_),
    .B1(_04713_),
    .B2(_04714_),
    .C1(_13384_),
    .Y(_04715_));
 sky130_fd_sc_hd__nand4_1 _15204_ (.A(_13364_),
    .B(_13371_),
    .C(_13378_),
    .D(_13385_),
    .Y(_04716_));
 sky130_fd_sc_hd__nor2_1 _15205_ (.A(_04660_),
    .B(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__and3_4 _15206_ (.A(_13357_),
    .B(_04678_),
    .C(_04717_),
    .X(_04718_));
 sky130_fd_sc_hd__o2111ai_1 _15207_ (.A1(_13300_),
    .A2(_04627_),
    .B1(_04650_),
    .C1(_04718_),
    .D1(_13308_),
    .Y(_04719_));
 sky130_fd_sc_hd__a21oi_1 _15208_ (.A1(_13315_),
    .A2(_13307_),
    .B1(_13314_),
    .Y(_04720_));
 sky130_fd_sc_hd__nor2_1 _15209_ (.A(_04641_),
    .B(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__o31ai_1 _15210_ (.A1(_13321_),
    .A2(_13328_),
    .A3(_04721_),
    .B1(_04718_),
    .Y(_04722_));
 sky130_fd_sc_hd__and3_4 _15211_ (.A(_04715_),
    .B(_04719_),
    .C(_04722_),
    .X(_04723_));
 sky130_fd_sc_hd__xnor2_2 _15212_ (.A(_13392_),
    .B(_04723_),
    .Y(_13393_));
 sky130_fd_sc_hd__inv_4 _15213_ (.A(_13393_),
    .Y(_12291_));
 sky130_fd_sc_hd__xnor2_1 _15214_ (.A(_04437_),
    .B(_04487_),
    .Y(_04724_));
 sky130_fd_sc_hd__xnor2_1 _15215_ (.A(_04499_),
    .B(_04724_),
    .Y(_12290_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1409 ();
 sky130_fd_sc_hd__xnor2_2 _15217_ (.A(_12968_),
    .B(_04480_),
    .Y(_04726_));
 sky130_fd_sc_hd__nand2_2 _15218_ (.A(\hash.CA2.a_dash[24] ),
    .B(_04726_),
    .Y(_04727_));
 sky130_fd_sc_hd__o21ai_0 _15219_ (.A1(\hash.CA2.a_dash[24] ),
    .A2(_04726_),
    .B1(\hash.CA2.b_dash[24] ),
    .Y(_04728_));
 sky130_fd_sc_hd__nand2_2 _15220_ (.A(_04727_),
    .B(_04728_),
    .Y(_04729_));
 sky130_fd_sc_hd__inv_4 _15221_ (.A(_04729_),
    .Y(_12301_));
 sky130_fd_sc_hd__a21o_1 _15222_ (.A1(_13385_),
    .A2(_04710_),
    .B1(_13384_),
    .X(_04730_));
 sky130_fd_sc_hd__a21oi_1 _15223_ (.A1(_13392_),
    .A2(_04730_),
    .B1(_13391_),
    .Y(_04731_));
 sky130_fd_sc_hd__xnor2_1 _15224_ (.A(_13399_),
    .B(_04731_),
    .Y(_13400_));
 sky130_fd_sc_hd__clkinv_2 _15225_ (.A(_13400_),
    .Y(_12300_));
 sky130_fd_sc_hd__xnor2_1 _15226_ (.A(_04475_),
    .B(_04501_),
    .Y(_04732_));
 sky130_fd_sc_hd__xnor2_1 _15227_ (.A(_04517_),
    .B(_04732_),
    .Y(_12299_));
 sky130_fd_sc_hd__inv_12 _15228_ (.A(\hash.CA2.b_dash[25] ),
    .Y(_04733_));
 sky130_fd_sc_hd__inv_4 _15229_ (.A(\hash.CA2.a_dash[25] ),
    .Y(_04734_));
 sky130_fd_sc_hd__maj3_1 _15230_ (.A(_04733_),
    .B(_04734_),
    .C(_04499_),
    .X(_12310_));
 sky130_fd_sc_hd__a21o_4 _15231_ (.A1(_13399_),
    .A2(_13391_),
    .B1(_13398_),
    .X(_04735_));
 sky130_fd_sc_hd__nand2_2 _15232_ (.A(_13392_),
    .B(_13399_),
    .Y(_04736_));
 sky130_fd_sc_hd__nor2_1 _15233_ (.A(_04723_),
    .B(_04736_),
    .Y(_04737_));
 sky130_fd_sc_hd__nor2_1 _15234_ (.A(_04735_),
    .B(_04737_),
    .Y(_04738_));
 sky130_fd_sc_hd__xnor2_1 _15235_ (.A(_13406_),
    .B(_04738_),
    .Y(_13407_));
 sky130_fd_sc_hd__inv_4 _15236_ (.A(_13407_),
    .Y(_12309_));
 sky130_fd_sc_hd__xor2_1 _15237_ (.A(_04484_),
    .B(_04522_),
    .X(_04739_));
 sky130_fd_sc_hd__xnor2_1 _15238_ (.A(net1073),
    .B(_04739_),
    .Y(_12308_));
 sky130_fd_sc_hd__maj3_2 _15239_ (.A(\hash.CA2.b_dash[26] ),
    .B(\hash.CA2.a_dash[26] ),
    .C(net1101),
    .X(_04740_));
 sky130_fd_sc_hd__inv_2 _15240_ (.A(_04740_),
    .Y(_12319_));
 sky130_fd_sc_hd__nand2_1 _15241_ (.A(_13385_),
    .B(_13406_),
    .Y(_04741_));
 sky130_fd_sc_hd__nor2_1 _15242_ (.A(_04736_),
    .B(_04741_),
    .Y(_04742_));
 sky130_fd_sc_hd__nand2_1 _15243_ (.A(_13406_),
    .B(_13384_),
    .Y(_04743_));
 sky130_fd_sc_hd__nand2_1 _15244_ (.A(_13406_),
    .B(_04735_),
    .Y(_04744_));
 sky130_fd_sc_hd__o21ai_0 _15245_ (.A1(_04736_),
    .A2(_04743_),
    .B1(_04744_),
    .Y(_04745_));
 sky130_fd_sc_hd__a211o_4 _15246_ (.A1(_04710_),
    .A2(_04742_),
    .B1(_04745_),
    .C1(_13405_),
    .X(_04746_));
 sky130_fd_sc_hd__xor2_4 _15247_ (.A(_13413_),
    .B(_04746_),
    .X(_13414_));
 sky130_fd_sc_hd__inv_4 _15248_ (.A(net1064),
    .Y(_12318_));
 sky130_fd_sc_hd__xnor2_1 _15249_ (.A(_04503_),
    .B(_04542_),
    .Y(_04747_));
 sky130_fd_sc_hd__xnor2_1 _15250_ (.A(_04662_),
    .B(_04747_),
    .Y(_12317_));
 sky130_fd_sc_hd__maj3_1 _15251_ (.A(\hash.CA2.b_dash[27] ),
    .B(\hash.CA2.a_dash[27] ),
    .C(_04537_),
    .X(_04748_));
 sky130_fd_sc_hd__inv_1 _15252_ (.A(_04748_),
    .Y(_12328_));
 sky130_fd_sc_hd__nand4_1 _15253_ (.A(_13392_),
    .B(_13399_),
    .C(_13406_),
    .D(_13413_),
    .Y(_04749_));
 sky130_fd_sc_hd__clkinv_1 _15254_ (.A(_04744_),
    .Y(_04750_));
 sky130_fd_sc_hd__o21ai_1 _15255_ (.A1(_13405_),
    .A2(_04750_),
    .B1(_13413_),
    .Y(_04751_));
 sky130_fd_sc_hd__o21ai_2 _15256_ (.A1(_04723_),
    .A2(_04749_),
    .B1(_04751_),
    .Y(_04752_));
 sky130_fd_sc_hd__nor2_4 _15257_ (.A(_13412_),
    .B(_04752_),
    .Y(_04753_));
 sky130_fd_sc_hd__xnor2_4 _15258_ (.A(_13420_),
    .B(_04753_),
    .Y(_13421_));
 sky130_fd_sc_hd__inv_1 _15259_ (.A(_13421_),
    .Y(_12327_));
 sky130_fd_sc_hd__a21oi_4 _15260_ (.A1(_04569_),
    .A2(_04570_),
    .B1(_04573_),
    .Y(_04754_));
 sky130_fd_sc_hd__xor2_1 _15261_ (.A(_04520_),
    .B(_04562_),
    .X(_04755_));
 sky130_fd_sc_hd__xnor2_1 _15262_ (.A(_04754_),
    .B(_04755_),
    .Y(_12326_));
 sky130_fd_sc_hd__nand2_2 _15263_ (.A(\hash.CA2.a_dash[28] ),
    .B(_04554_),
    .Y(_04756_));
 sky130_fd_sc_hd__o21ai_0 _15264_ (.A1(\hash.CA2.a_dash[28] ),
    .A2(_04554_),
    .B1(\hash.CA2.b_dash[28] ),
    .Y(_04757_));
 sky130_fd_sc_hd__nand2_1 _15265_ (.A(_04756_),
    .B(_04757_),
    .Y(_04758_));
 sky130_fd_sc_hd__inv_2 _15266_ (.A(_04758_),
    .Y(_12337_));
 sky130_fd_sc_hd__a21o_1 _15267_ (.A1(_13413_),
    .A2(_04746_),
    .B1(_13412_),
    .X(_04759_));
 sky130_fd_sc_hd__a21oi_2 _15268_ (.A1(_13420_),
    .A2(_04759_),
    .B1(_13419_),
    .Y(_04760_));
 sky130_fd_sc_hd__xor2_2 _15269_ (.A(_13427_),
    .B(_04760_),
    .X(_12336_));
 sky130_fd_sc_hd__xnor2_1 _15270_ (.A(_04541_),
    .B(_04580_),
    .Y(_04761_));
 sky130_fd_sc_hd__xnor2_1 _15271_ (.A(net1095),
    .B(_04761_),
    .Y(_12335_));
 sky130_fd_sc_hd__nor2_1 _15272_ (.A(\hash.CA2.a_dash[29] ),
    .B(_04754_),
    .Y(_04762_));
 sky130_fd_sc_hd__a21oi_1 _15273_ (.A1(\hash.CA2.a_dash[29] ),
    .A2(_04754_),
    .B1(\hash.CA2.b_dash[29] ),
    .Y(_04763_));
 sky130_fd_sc_hd__nor2_1 _15274_ (.A(_04762_),
    .B(_04763_),
    .Y(_04764_));
 sky130_fd_sc_hd__clkinvlp_2 _15275_ (.A(_04764_),
    .Y(_12346_));
 sky130_fd_sc_hd__inv_1 _15276_ (.A(_13420_),
    .Y(_04765_));
 sky130_fd_sc_hd__o21bai_1 _15277_ (.A1(_04765_),
    .A2(_04753_),
    .B1_N(_13419_),
    .Y(_04766_));
 sky130_fd_sc_hd__a21oi_1 _15278_ (.A1(_13427_),
    .A2(_04766_),
    .B1(_13426_),
    .Y(_04767_));
 sky130_fd_sc_hd__xnor2_2 _15279_ (.A(_13434_),
    .B(_04767_),
    .Y(_13435_));
 sky130_fd_sc_hd__inv_1 _15280_ (.A(_13435_),
    .Y(_12345_));
 sky130_fd_sc_hd__xor2_1 _15281_ (.A(_04559_),
    .B(_04599_),
    .X(_04768_));
 sky130_fd_sc_hd__xnor2_1 _15282_ (.A(_04612_),
    .B(_04768_),
    .Y(_12344_));
 sky130_fd_sc_hd__clkinvlp_4 _15283_ (.A(\hash.CA2.a_dash[30] ),
    .Y(_04769_));
 sky130_fd_sc_hd__nand2_2 _15284_ (.A(_04769_),
    .B(net1095),
    .Y(_04770_));
 sky130_fd_sc_hd__nor2_2 _15285_ (.A(_04769_),
    .B(net1095),
    .Y(_04771_));
 sky130_fd_sc_hd__a21oi_2 _15286_ (.A1(\hash.CA2.b_dash[30] ),
    .A2(_04770_),
    .B1(_04771_),
    .Y(_12355_));
 sky130_fd_sc_hd__nand2_1 _15287_ (.A(_13413_),
    .B(_04746_),
    .Y(_04772_));
 sky130_fd_sc_hd__a21oi_1 _15288_ (.A1(_13427_),
    .A2(_13419_),
    .B1(_13426_),
    .Y(_04773_));
 sky130_fd_sc_hd__nor2b_2 _15289_ (.A(_04773_),
    .B_N(_13434_),
    .Y(_04774_));
 sky130_fd_sc_hd__nor3_2 _15290_ (.A(_13412_),
    .B(_13433_),
    .C(_04774_),
    .Y(_04775_));
 sky130_fd_sc_hd__a311o_1 _15291_ (.A1(_13420_),
    .A2(_13427_),
    .A3(_13434_),
    .B1(_13433_),
    .C1(_04774_),
    .X(_04776_));
 sky130_fd_sc_hd__a21boi_2 _15292_ (.A1(_04772_),
    .A2(_04775_),
    .B1_N(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__xnor2_2 _15293_ (.A(_13441_),
    .B(_04777_),
    .Y(_12354_));
 sky130_fd_sc_hd__xnor2_1 _15294_ (.A(_12922_),
    .B(_04614_),
    .Y(_04778_));
 sky130_fd_sc_hd__xnor2_1 _15295_ (.A(_04681_),
    .B(_04778_),
    .Y(_12353_));
 sky130_fd_sc_hd__nor2_1 _15296_ (.A(net342),
    .B(_13445_),
    .Y(_00781_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1408 ();
 sky130_fd_sc_hd__or2_0 _15298_ (.A(net344),
    .B(net1121),
    .X(\hash.CA1.f[2] ));
 sky130_fd_sc_hd__inv_2 _15299_ (.A(\hash.CA1.f[2] ),
    .Y(_00813_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1404 ();
 sky130_fd_sc_hd__nor2_1 _15304_ (.A(net344),
    .B(\hash.CA2.S1.X[3] ),
    .Y(_13851_));
 sky130_fd_sc_hd__nor2b_4 _15305_ (.A(net1038),
    .B_N(_13528_),
    .Y(_04784_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1403 ();
 sky130_fd_sc_hd__nand2_8 _15307_ (.A(_09735_),
    .B(_04784_),
    .Y(_04786_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1400 ();
 sky130_fd_sc_hd__mux2i_4 _15311_ (.A0(_12986_),
    .A1(\w[62][0] ),
    .S(net353),
    .Y(_04790_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1398 ();
 sky130_fd_sc_hd__nand2_1 _15314_ (.A(net245),
    .B(_04786_),
    .Y(_04793_));
 sky130_fd_sc_hd__o21ai_0 _15315_ (.A1(_04786_),
    .A2(_04790_),
    .B1(_04793_),
    .Y(_00129_));
 sky130_fd_sc_hd__mux2i_4 _15316_ (.A0(_12989_),
    .A1(\w[62][1] ),
    .S(net352),
    .Y(_04794_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1397 ();
 sky130_fd_sc_hd__nand2_1 _15318_ (.A(net234),
    .B(_04786_),
    .Y(_04796_));
 sky130_fd_sc_hd__o21ai_0 _15319_ (.A1(_04786_),
    .A2(_04794_),
    .B1(_04796_),
    .Y(_00140_));
 sky130_fd_sc_hd__clkinv_16 _15320_ (.A(net356),
    .Y(_04797_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1395 ();
 sky130_fd_sc_hd__nand2_2 _15323_ (.A(_11602_),
    .B(_04797_),
    .Y(_04800_));
 sky130_fd_sc_hd__o21ai_4 _15324_ (.A1(\w[62][2] ),
    .A2(_04797_),
    .B1(_04800_),
    .Y(_04801_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1394 ();
 sky130_fd_sc_hd__nand2_1 _15326_ (.A(net222),
    .B(_04786_),
    .Y(_04803_));
 sky130_fd_sc_hd__o21ai_0 _15327_ (.A1(_04786_),
    .A2(_04801_),
    .B1(_04803_),
    .Y(_00151_));
 sky130_fd_sc_hd__nor2b_2 _15328_ (.A(_12997_),
    .B_N(_11601_),
    .Y(_04804_));
 sky130_fd_sc_hd__nor2b_4 _15329_ (.A(_11601_),
    .B_N(_12997_),
    .Y(_04805_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1393 ();
 sky130_fd_sc_hd__o21ai_4 _15331_ (.A1(_04804_),
    .A2(_04805_),
    .B1(_04797_),
    .Y(_04807_));
 sky130_fd_sc_hd__o21ai_4 _15332_ (.A1(\w[62][3] ),
    .A2(_04797_),
    .B1(_04807_),
    .Y(_04808_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1392 ();
 sky130_fd_sc_hd__nand2_1 _15334_ (.A(net211),
    .B(_04786_),
    .Y(_04810_));
 sky130_fd_sc_hd__o21ai_0 _15335_ (.A1(_04786_),
    .A2(_04808_),
    .B1(_04810_),
    .Y(_00154_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1391 ();
 sky130_fd_sc_hd__clkinv_1 _15337_ (.A(_13001_),
    .Y(_04812_));
 sky130_fd_sc_hd__a21o_1 _15338_ (.A1(_12988_),
    .A2(_12993_),
    .B1(_12992_),
    .X(_04813_));
 sky130_fd_sc_hd__a21oi_2 _15339_ (.A1(_12997_),
    .A2(_04813_),
    .B1(_12996_),
    .Y(_04814_));
 sky130_fd_sc_hd__xnor2_2 _15340_ (.A(_04812_),
    .B(_04814_),
    .Y(_04815_));
 sky130_fd_sc_hd__nand2_8 _15341_ (.A(_04797_),
    .B(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__o21ai_4 _15342_ (.A1(\w[62][4] ),
    .A2(_04797_),
    .B1(_04816_),
    .Y(_04817_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1390 ();
 sky130_fd_sc_hd__nand2_1 _15344_ (.A(net200),
    .B(_04786_),
    .Y(_04819_));
 sky130_fd_sc_hd__o21ai_0 _15345_ (.A1(_04786_),
    .A2(_04817_),
    .B1(_04819_),
    .Y(_00155_));
 sky130_fd_sc_hd__inv_2 _15346_ (.A(_13000_),
    .Y(_04820_));
 sky130_fd_sc_hd__o21ai_2 _15347_ (.A1(_12996_),
    .A2(_04805_),
    .B1(_13001_),
    .Y(_04821_));
 sky130_fd_sc_hd__a21boi_4 _15348_ (.A1(_04820_),
    .A2(_04821_),
    .B1_N(_13005_),
    .Y(_04822_));
 sky130_fd_sc_hd__nand2_1 _15349_ (.A(_04820_),
    .B(_04821_),
    .Y(_04823_));
 sky130_fd_sc_hd__nor2_1 _15350_ (.A(_13005_),
    .B(_04823_),
    .Y(_04824_));
 sky130_fd_sc_hd__o21ai_4 _15351_ (.A1(_04822_),
    .A2(_04824_),
    .B1(_04797_),
    .Y(_04825_));
 sky130_fd_sc_hd__o21ai_4 _15352_ (.A1(\w[62][5] ),
    .A2(_04797_),
    .B1(_04825_),
    .Y(_04826_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1389 ();
 sky130_fd_sc_hd__nand2_1 _15354_ (.A(net189),
    .B(_04786_),
    .Y(_04828_));
 sky130_fd_sc_hd__o21ai_0 _15355_ (.A1(_04786_),
    .A2(_04826_),
    .B1(_04828_),
    .Y(_00156_));
 sky130_fd_sc_hd__inv_2 _15356_ (.A(_13009_),
    .Y(_04829_));
 sky130_fd_sc_hd__o21ai_0 _15357_ (.A1(_04812_),
    .A2(_04814_),
    .B1(_04820_),
    .Y(_04830_));
 sky130_fd_sc_hd__a21oi_2 _15358_ (.A1(_13005_),
    .A2(_04830_),
    .B1(_13004_),
    .Y(_04831_));
 sky130_fd_sc_hd__xnor2_1 _15359_ (.A(_04829_),
    .B(_04831_),
    .Y(_04832_));
 sky130_fd_sc_hd__nand2_2 _15360_ (.A(_04797_),
    .B(_04832_),
    .Y(_04833_));
 sky130_fd_sc_hd__o21ai_4 _15361_ (.A1(\w[62][6] ),
    .A2(_04797_),
    .B1(_04833_),
    .Y(_04834_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1388 ();
 sky130_fd_sc_hd__nand2_1 _15363_ (.A(net178),
    .B(_04786_),
    .Y(_04836_));
 sky130_fd_sc_hd__o21ai_0 _15364_ (.A1(_04786_),
    .A2(_04834_),
    .B1(_04836_),
    .Y(_00157_));
 sky130_fd_sc_hd__clkinv_4 _15365_ (.A(_13008_),
    .Y(_04837_));
 sky130_fd_sc_hd__o21ai_2 _15366_ (.A1(_13004_),
    .A2(_04822_),
    .B1(_13009_),
    .Y(_04838_));
 sky130_fd_sc_hd__a21boi_4 _15367_ (.A1(_04837_),
    .A2(_04838_),
    .B1_N(_13013_),
    .Y(_04839_));
 sky130_fd_sc_hd__nand2_1 _15368_ (.A(_04837_),
    .B(_04838_),
    .Y(_04840_));
 sky130_fd_sc_hd__nor2_1 _15369_ (.A(_13013_),
    .B(_04840_),
    .Y(_04841_));
 sky130_fd_sc_hd__o21ai_4 _15370_ (.A1(_04839_),
    .A2(_04841_),
    .B1(_04797_),
    .Y(_04842_));
 sky130_fd_sc_hd__o21ai_4 _15371_ (.A1(\w[62][7] ),
    .A2(_04797_),
    .B1(_04842_),
    .Y(_04843_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1387 ();
 sky130_fd_sc_hd__nand2_1 _15373_ (.A(net167),
    .B(_04786_),
    .Y(_04845_));
 sky130_fd_sc_hd__o21ai_0 _15374_ (.A1(_04786_),
    .A2(_04843_),
    .B1(_04845_),
    .Y(_00158_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1385 ();
 sky130_fd_sc_hd__o21ai_4 _15377_ (.A1(_04829_),
    .A2(_04831_),
    .B1(_04837_),
    .Y(_04848_));
 sky130_fd_sc_hd__a21oi_2 _15378_ (.A1(_13013_),
    .A2(_04848_),
    .B1(_13012_),
    .Y(_04849_));
 sky130_fd_sc_hd__xor2_2 _15379_ (.A(_13017_),
    .B(_04849_),
    .X(_04850_));
 sky130_fd_sc_hd__nor2_1 _15380_ (.A(net354),
    .B(_04850_),
    .Y(_04851_));
 sky130_fd_sc_hd__a21oi_4 _15381_ (.A1(\w[62][8] ),
    .A2(net354),
    .B1(_04851_),
    .Y(_04852_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1384 ();
 sky130_fd_sc_hd__nand2_1 _15383_ (.A(net156),
    .B(_04786_),
    .Y(_04854_));
 sky130_fd_sc_hd__o21ai_0 _15384_ (.A1(_04786_),
    .A2(_04852_),
    .B1(_04854_),
    .Y(_00159_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1383 ();
 sky130_fd_sc_hd__o21ai_0 _15386_ (.A1(_13012_),
    .A2(_04839_),
    .B1(_13017_),
    .Y(_04856_));
 sky130_fd_sc_hd__nand2b_1 _15387_ (.A_N(_13016_),
    .B(_04856_),
    .Y(_04857_));
 sky130_fd_sc_hd__xnor2_1 _15388_ (.A(_13021_),
    .B(_04857_),
    .Y(_04858_));
 sky130_fd_sc_hd__nor2_4 _15389_ (.A(net352),
    .B(_04858_),
    .Y(_04859_));
 sky130_fd_sc_hd__a21oi_4 _15390_ (.A1(\w[62][9] ),
    .A2(net354),
    .B1(_04859_),
    .Y(_04860_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1382 ();
 sky130_fd_sc_hd__nand2_1 _15392_ (.A(net145),
    .B(_04786_),
    .Y(_04862_));
 sky130_fd_sc_hd__o21ai_0 _15393_ (.A1(_04786_),
    .A2(_04860_),
    .B1(_04862_),
    .Y(_00160_));
 sky130_fd_sc_hd__clkinv_1 _15394_ (.A(_13020_),
    .Y(_04863_));
 sky130_fd_sc_hd__a211o_4 _15395_ (.A1(_13013_),
    .A2(_04848_),
    .B1(_13016_),
    .C1(_13012_),
    .X(_04864_));
 sky130_fd_sc_hd__o21a_4 _15396_ (.A1(_13017_),
    .A2(_13016_),
    .B1(_13021_),
    .X(_04865_));
 sky130_fd_sc_hd__nand2_1 _15397_ (.A(_04864_),
    .B(_04865_),
    .Y(_04866_));
 sky130_fd_sc_hd__inv_1 _15398_ (.A(_13025_),
    .Y(_04867_));
 sky130_fd_sc_hd__a21oi_2 _15399_ (.A1(_04863_),
    .A2(_04866_),
    .B1(_04867_),
    .Y(_04868_));
 sky130_fd_sc_hd__and3_4 _15400_ (.A(_04867_),
    .B(_04863_),
    .C(_04866_),
    .X(_04869_));
 sky130_fd_sc_hd__nor3_4 _15401_ (.A(net352),
    .B(_04868_),
    .C(_04869_),
    .Y(_04870_));
 sky130_fd_sc_hd__a21oi_4 _15402_ (.A1(\w[62][10] ),
    .A2(net354),
    .B1(_04870_),
    .Y(_04871_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1380 ();
 sky130_fd_sc_hd__nand2_1 _15405_ (.A(net134),
    .B(_04786_),
    .Y(_04874_));
 sky130_fd_sc_hd__o21ai_0 _15406_ (.A1(_04786_),
    .A2(_04871_),
    .B1(_04874_),
    .Y(_00130_));
 sky130_fd_sc_hd__nand2_1 _15407_ (.A(_13021_),
    .B(_13016_),
    .Y(_04875_));
 sky130_fd_sc_hd__nand2_1 _15408_ (.A(_04863_),
    .B(_04875_),
    .Y(_04876_));
 sky130_fd_sc_hd__a21oi_2 _15409_ (.A1(_13025_),
    .A2(_04876_),
    .B1(_13024_),
    .Y(_04877_));
 sky130_fd_sc_hd__o2111ai_2 _15410_ (.A1(_13012_),
    .A2(_04839_),
    .B1(_13017_),
    .C1(_13021_),
    .D1(_13025_),
    .Y(_04878_));
 sky130_fd_sc_hd__a21boi_4 _15411_ (.A1(_04877_),
    .A2(_04878_),
    .B1_N(_13029_),
    .Y(_04879_));
 sky130_fd_sc_hd__nand2_1 _15412_ (.A(_04877_),
    .B(_04878_),
    .Y(_04880_));
 sky130_fd_sc_hd__nor2_1 _15413_ (.A(_13029_),
    .B(_04880_),
    .Y(_04881_));
 sky130_fd_sc_hd__o21ai_2 _15414_ (.A1(_04879_),
    .A2(_04881_),
    .B1(_04797_),
    .Y(_04882_));
 sky130_fd_sc_hd__o21ai_4 _15415_ (.A1(\w[62][11] ),
    .A2(_04797_),
    .B1(_04882_),
    .Y(_04883_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1379 ();
 sky130_fd_sc_hd__nand2_1 _15417_ (.A(net123),
    .B(_04786_),
    .Y(_04885_));
 sky130_fd_sc_hd__o21ai_0 _15418_ (.A1(_04786_),
    .A2(_04883_),
    .B1(_04885_),
    .Y(_00131_));
 sky130_fd_sc_hd__a2111oi_4 _15419_ (.A1(_04864_),
    .A2(_04865_),
    .B1(_13020_),
    .C1(_13024_),
    .D1(_13028_),
    .Y(_04886_));
 sky130_fd_sc_hd__or2_4 _15420_ (.A(_13025_),
    .B(_13024_),
    .X(_04887_));
 sky130_fd_sc_hd__a21oi_4 _15421_ (.A1(_13029_),
    .A2(_04887_),
    .B1(_13028_),
    .Y(_04888_));
 sky130_fd_sc_hd__nor2_4 _15422_ (.A(_04886_),
    .B(_04888_),
    .Y(_04889_));
 sky130_fd_sc_hd__xnor2_2 _15423_ (.A(_13033_),
    .B(_04889_),
    .Y(_04890_));
 sky130_fd_sc_hd__nand2_2 _15424_ (.A(_04797_),
    .B(_04890_),
    .Y(_04891_));
 sky130_fd_sc_hd__o21ai_4 _15425_ (.A1(\w[62][12] ),
    .A2(_04797_),
    .B1(_04891_),
    .Y(_04892_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1378 ();
 sky130_fd_sc_hd__nand2_1 _15427_ (.A(net111),
    .B(_04786_),
    .Y(_04894_));
 sky130_fd_sc_hd__o21ai_0 _15428_ (.A1(_04786_),
    .A2(_04892_),
    .B1(_04894_),
    .Y(_00132_));
 sky130_fd_sc_hd__or2_4 _15429_ (.A(_13028_),
    .B(_04879_),
    .X(_04895_));
 sky130_fd_sc_hd__a21o_1 _15430_ (.A1(_13033_),
    .A2(_04895_),
    .B1(_13032_),
    .X(_04896_));
 sky130_fd_sc_hd__xnor2_1 _15431_ (.A(_13037_),
    .B(_04896_),
    .Y(_04897_));
 sky130_fd_sc_hd__nand2_2 _15432_ (.A(_04797_),
    .B(_04897_),
    .Y(_04898_));
 sky130_fd_sc_hd__o21ai_4 _15433_ (.A1(\w[62][13] ),
    .A2(_04797_),
    .B1(_04898_),
    .Y(_04899_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1377 ();
 sky130_fd_sc_hd__nand2_1 _15435_ (.A(net100),
    .B(_04786_),
    .Y(_04901_));
 sky130_fd_sc_hd__o21ai_0 _15436_ (.A1(_04786_),
    .A2(_04899_),
    .B1(_04901_),
    .Y(_00133_));
 sky130_fd_sc_hd__a21o_1 _15437_ (.A1(_13033_),
    .A2(_04889_),
    .B1(_13032_),
    .X(_04902_));
 sky130_fd_sc_hd__a21oi_1 _15438_ (.A1(_13037_),
    .A2(_04902_),
    .B1(_13036_),
    .Y(_04903_));
 sky130_fd_sc_hd__xor2_1 _15439_ (.A(_13041_),
    .B(_04903_),
    .X(_04904_));
 sky130_fd_sc_hd__nor2_2 _15440_ (.A(net354),
    .B(_04904_),
    .Y(_04905_));
 sky130_fd_sc_hd__a21oi_4 _15441_ (.A1(\w[62][14] ),
    .A2(net354),
    .B1(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1376 ();
 sky130_fd_sc_hd__nand2_1 _15443_ (.A(net89),
    .B(_04786_),
    .Y(_04908_));
 sky130_fd_sc_hd__o21ai_0 _15444_ (.A1(_04786_),
    .A2(_04906_),
    .B1(_04908_),
    .Y(_00134_));
 sky130_fd_sc_hd__a21o_1 _15445_ (.A1(_13037_),
    .A2(_04896_),
    .B1(_13036_),
    .X(_04909_));
 sky130_fd_sc_hd__a21oi_2 _15446_ (.A1(_13041_),
    .A2(_04909_),
    .B1(_13040_),
    .Y(_04910_));
 sky130_fd_sc_hd__xnor2_4 _15447_ (.A(_13045_),
    .B(_04910_),
    .Y(_04911_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1375 ();
 sky130_fd_sc_hd__mux2i_4 _15449_ (.A0(\w[62][15] ),
    .A1(_04911_),
    .S(_04797_),
    .Y(_04913_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1374 ();
 sky130_fd_sc_hd__nand2_1 _15451_ (.A(net78),
    .B(_04786_),
    .Y(_04915_));
 sky130_fd_sc_hd__o21ai_0 _15452_ (.A1(_04786_),
    .A2(_04913_),
    .B1(_04915_),
    .Y(_00135_));
 sky130_fd_sc_hd__nand4_1 _15453_ (.A(_13033_),
    .B(_13037_),
    .C(_13041_),
    .D(_13045_),
    .Y(_04916_));
 sky130_fd_sc_hd__a21o_1 _15454_ (.A1(_13037_),
    .A2(_13032_),
    .B1(_13036_),
    .X(_04917_));
 sky130_fd_sc_hd__a21o_1 _15455_ (.A1(_13041_),
    .A2(_04917_),
    .B1(_13040_),
    .X(_04918_));
 sky130_fd_sc_hd__a21oi_2 _15456_ (.A1(_13045_),
    .A2(_04918_),
    .B1(_13044_),
    .Y(_04919_));
 sky130_fd_sc_hd__o31ai_1 _15457_ (.A1(_04886_),
    .A2(_04888_),
    .A3(_04916_),
    .B1(_04919_),
    .Y(_04920_));
 sky130_fd_sc_hd__xnor2_1 _15458_ (.A(_13049_),
    .B(_04920_),
    .Y(_04921_));
 sky130_fd_sc_hd__nand2_2 _15459_ (.A(_04797_),
    .B(_04921_),
    .Y(_04922_));
 sky130_fd_sc_hd__o21ai_4 _15460_ (.A1(\w[62][16] ),
    .A2(_04797_),
    .B1(_04922_),
    .Y(_04923_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1373 ();
 sky130_fd_sc_hd__nand2_1 _15462_ (.A(net67),
    .B(_04786_),
    .Y(_04925_));
 sky130_fd_sc_hd__o21ai_0 _15463_ (.A1(_04786_),
    .A2(_04923_),
    .B1(_04925_),
    .Y(_00136_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1372 ();
 sky130_fd_sc_hd__nor2_1 _15465_ (.A(_13028_),
    .B(_04879_),
    .Y(_04927_));
 sky130_fd_sc_hd__o21ai_0 _15466_ (.A1(_04927_),
    .A2(_04916_),
    .B1(_04919_),
    .Y(_04928_));
 sky130_fd_sc_hd__a21oi_1 _15467_ (.A1(_13049_),
    .A2(_04928_),
    .B1(_13048_),
    .Y(_04929_));
 sky130_fd_sc_hd__xor2_2 _15468_ (.A(_13053_),
    .B(_04929_),
    .X(_04930_));
 sky130_fd_sc_hd__nor2_2 _15469_ (.A(net353),
    .B(_04930_),
    .Y(_04931_));
 sky130_fd_sc_hd__a21oi_4 _15470_ (.A1(\w[62][17] ),
    .A2(net353),
    .B1(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1371 ();
 sky130_fd_sc_hd__nand2_1 _15472_ (.A(net56),
    .B(_04786_),
    .Y(_04934_));
 sky130_fd_sc_hd__o21ai_0 _15473_ (.A1(_04786_),
    .A2(_04932_),
    .B1(_04934_),
    .Y(_00137_));
 sky130_fd_sc_hd__a21o_1 _15474_ (.A1(_13049_),
    .A2(_04920_),
    .B1(_13048_),
    .X(_04935_));
 sky130_fd_sc_hd__a21oi_1 _15475_ (.A1(_13053_),
    .A2(_04935_),
    .B1(_13052_),
    .Y(_04936_));
 sky130_fd_sc_hd__xor2_1 _15476_ (.A(_13057_),
    .B(_04936_),
    .X(_04937_));
 sky130_fd_sc_hd__nor2_1 _15477_ (.A(net352),
    .B(_04937_),
    .Y(_04938_));
 sky130_fd_sc_hd__a21oi_4 _15478_ (.A1(\w[62][18] ),
    .A2(net352),
    .B1(_04938_),
    .Y(_04939_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1370 ();
 sky130_fd_sc_hd__nand2_1 _15480_ (.A(net45),
    .B(_04786_),
    .Y(_04941_));
 sky130_fd_sc_hd__o21ai_0 _15481_ (.A1(_04786_),
    .A2(_04939_),
    .B1(_04941_),
    .Y(_00138_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1369 ();
 sky130_fd_sc_hd__nand3_1 _15483_ (.A(_13049_),
    .B(_13053_),
    .C(_13057_),
    .Y(_04943_));
 sky130_fd_sc_hd__nor2_2 _15484_ (.A(_04916_),
    .B(_04943_),
    .Y(_04944_));
 sky130_fd_sc_hd__a21o_1 _15485_ (.A1(_13053_),
    .A2(_13048_),
    .B1(_13052_),
    .X(_04945_));
 sky130_fd_sc_hd__a21o_4 _15486_ (.A1(_13057_),
    .A2(_04945_),
    .B1(_13056_),
    .X(_04946_));
 sky130_fd_sc_hd__or2_4 _15487_ (.A(_04919_),
    .B(_04943_),
    .X(_04947_));
 sky130_fd_sc_hd__nand2b_2 _15488_ (.A_N(_04946_),
    .B(_04947_),
    .Y(_04948_));
 sky130_fd_sc_hd__a21oi_2 _15489_ (.A1(_04895_),
    .A2(_04944_),
    .B1(_04948_),
    .Y(_04949_));
 sky130_fd_sc_hd__xnor2_2 _15490_ (.A(_13061_),
    .B(_04949_),
    .Y(_04950_));
 sky130_fd_sc_hd__mux2i_4 _15491_ (.A0(\w[62][19] ),
    .A1(_04950_),
    .S(_04797_),
    .Y(_04951_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1368 ();
 sky130_fd_sc_hd__nand2_1 _15493_ (.A(net34),
    .B(_04786_),
    .Y(_04953_));
 sky130_fd_sc_hd__o21ai_0 _15494_ (.A1(_04786_),
    .A2(_04951_),
    .B1(_04953_),
    .Y(_00139_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1367 ();
 sky130_fd_sc_hd__a21oi_1 _15496_ (.A1(_13061_),
    .A2(_04948_),
    .B1(_13060_),
    .Y(_04955_));
 sky130_fd_sc_hd__inv_1 _15497_ (.A(_04955_),
    .Y(_04956_));
 sky130_fd_sc_hd__a31oi_1 _15498_ (.A1(_13061_),
    .A2(_04889_),
    .A3(_04944_),
    .B1(_04956_),
    .Y(_04957_));
 sky130_fd_sc_hd__xor2_1 _15499_ (.A(_13065_),
    .B(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__nor2_2 _15500_ (.A(net352),
    .B(_04958_),
    .Y(_04959_));
 sky130_fd_sc_hd__a21oi_4 _15501_ (.A1(\w[62][20] ),
    .A2(net352),
    .B1(_04959_),
    .Y(_04960_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1365 ();
 sky130_fd_sc_hd__nand2_1 _15504_ (.A(net23),
    .B(_04786_),
    .Y(_04963_));
 sky130_fd_sc_hd__o21ai_0 _15505_ (.A1(_04786_),
    .A2(_04960_),
    .B1(_04963_),
    .Y(_00141_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1364 ();
 sky130_fd_sc_hd__nand4_1 _15507_ (.A(_13049_),
    .B(_13053_),
    .C(_13057_),
    .D(_13028_),
    .Y(_04965_));
 sky130_fd_sc_hd__o21ai_0 _15508_ (.A1(_04916_),
    .A2(_04965_),
    .B1(_04947_),
    .Y(_04966_));
 sky130_fd_sc_hd__a21oi_2 _15509_ (.A1(_04879_),
    .A2(_04944_),
    .B1(_04966_),
    .Y(_04967_));
 sky130_fd_sc_hd__nor3_2 _15510_ (.A(_13060_),
    .B(_13064_),
    .C(_04946_),
    .Y(_04968_));
 sky130_fd_sc_hd__or2_0 _15511_ (.A(_13061_),
    .B(_13060_),
    .X(_04969_));
 sky130_fd_sc_hd__a21oi_2 _15512_ (.A1(_13065_),
    .A2(_04969_),
    .B1(_13064_),
    .Y(_04970_));
 sky130_fd_sc_hd__a21oi_2 _15513_ (.A1(_04967_),
    .A2(_04968_),
    .B1(_04970_),
    .Y(_04971_));
 sky130_fd_sc_hd__xnor2_1 _15514_ (.A(_13069_),
    .B(_04971_),
    .Y(_04972_));
 sky130_fd_sc_hd__nand2_2 _15515_ (.A(_04797_),
    .B(_04972_),
    .Y(_04973_));
 sky130_fd_sc_hd__o21ai_4 _15516_ (.A1(\w[62][21] ),
    .A2(_04797_),
    .B1(_04973_),
    .Y(_04974_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1363 ();
 sky130_fd_sc_hd__nand2_1 _15518_ (.A(net12),
    .B(_04786_),
    .Y(_04976_));
 sky130_fd_sc_hd__o21ai_0 _15519_ (.A1(_04786_),
    .A2(_04974_),
    .B1(_04976_),
    .Y(_00142_));
 sky130_fd_sc_hd__nand3_1 _15520_ (.A(_13061_),
    .B(_13065_),
    .C(_04944_),
    .Y(_04977_));
 sky130_fd_sc_hd__nor3_2 _15521_ (.A(_04886_),
    .B(_04888_),
    .C(_04977_),
    .Y(_04978_));
 sky130_fd_sc_hd__nor2b_2 _15522_ (.A(_04955_),
    .B_N(_13065_),
    .Y(_04979_));
 sky130_fd_sc_hd__o31ai_1 _15523_ (.A1(_13064_),
    .A2(_04978_),
    .A3(_04979_),
    .B1(_13069_),
    .Y(_04980_));
 sky130_fd_sc_hd__nand2b_2 _15524_ (.A_N(_13068_),
    .B(_04980_),
    .Y(_04981_));
 sky130_fd_sc_hd__xnor2_2 _15525_ (.A(_13073_),
    .B(_04981_),
    .Y(_04982_));
 sky130_fd_sc_hd__nor2_4 _15526_ (.A(net353),
    .B(_04982_),
    .Y(_04983_));
 sky130_fd_sc_hd__a21oi_4 _15527_ (.A1(\w[62][22] ),
    .A2(net353),
    .B1(_04983_),
    .Y(_04984_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1362 ();
 sky130_fd_sc_hd__nand2_1 _15529_ (.A(net779),
    .B(_04786_),
    .Y(_04986_));
 sky130_fd_sc_hd__o21ai_0 _15530_ (.A1(_04786_),
    .A2(_04984_),
    .B1(_04986_),
    .Y(_00143_));
 sky130_fd_sc_hd__a21o_1 _15531_ (.A1(_13069_),
    .A2(_04971_),
    .B1(_13068_),
    .X(_04987_));
 sky130_fd_sc_hd__a21oi_2 _15532_ (.A1(_13073_),
    .A2(_04987_),
    .B1(_13072_),
    .Y(_04988_));
 sky130_fd_sc_hd__xnor2_4 _15533_ (.A(_13077_),
    .B(_04988_),
    .Y(_04989_));
 sky130_fd_sc_hd__mux2i_4 _15534_ (.A0(\w[62][23] ),
    .A1(_04989_),
    .S(_04797_),
    .Y(_04990_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1361 ();
 sky130_fd_sc_hd__nand2_1 _15536_ (.A(net768),
    .B(_04786_),
    .Y(_04992_));
 sky130_fd_sc_hd__o21ai_0 _15537_ (.A1(_04786_),
    .A2(_04990_),
    .B1(_04992_),
    .Y(_00144_));
 sky130_fd_sc_hd__and3_1 _15538_ (.A(_13069_),
    .B(_13073_),
    .C(_13077_),
    .X(_04993_));
 sky130_fd_sc_hd__o31ai_2 _15539_ (.A1(_13064_),
    .A2(_04978_),
    .A3(_04979_),
    .B1(_04993_),
    .Y(_04994_));
 sky130_fd_sc_hd__and2_4 _15540_ (.A(_13073_),
    .B(_13068_),
    .X(_04995_));
 sky130_fd_sc_hd__o21ai_2 _15541_ (.A1(_13072_),
    .A2(_04995_),
    .B1(_13077_),
    .Y(_04996_));
 sky130_fd_sc_hd__nand3b_1 _15542_ (.A_N(_13076_),
    .B(_04994_),
    .C(_04996_),
    .Y(_04997_));
 sky130_fd_sc_hd__xnor2_2 _15543_ (.A(_13081_),
    .B(_04997_),
    .Y(_04998_));
 sky130_fd_sc_hd__nor2_2 _15544_ (.A(net353),
    .B(_04998_),
    .Y(_04999_));
 sky130_fd_sc_hd__a21oi_4 _15545_ (.A1(\w[62][24] ),
    .A2(net353),
    .B1(_04999_),
    .Y(_05000_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1360 ();
 sky130_fd_sc_hd__nand2_1 _15547_ (.A(net757),
    .B(_04786_),
    .Y(_05002_));
 sky130_fd_sc_hd__o21ai_0 _15548_ (.A1(_04786_),
    .A2(net1129),
    .B1(_05002_),
    .Y(_00145_));
 sky130_fd_sc_hd__nand4_1 _15549_ (.A(_13069_),
    .B(_13073_),
    .C(_13077_),
    .D(_13081_),
    .Y(_05003_));
 sky130_fd_sc_hd__a211oi_4 _15550_ (.A1(_04967_),
    .A2(_04968_),
    .B1(_04970_),
    .C1(_05003_),
    .Y(_05004_));
 sky130_fd_sc_hd__o211a_4 _15551_ (.A1(_13072_),
    .A2(_04995_),
    .B1(_13077_),
    .C1(_13081_),
    .X(_05005_));
 sky130_fd_sc_hd__nor2_4 _15552_ (.A(_05004_),
    .B(_05005_),
    .Y(_05006_));
 sky130_fd_sc_hd__a21oi_1 _15553_ (.A1(_13081_),
    .A2(_13076_),
    .B1(_13080_),
    .Y(_05007_));
 sky130_fd_sc_hd__nand2_1 _15554_ (.A(_05006_),
    .B(_05007_),
    .Y(_05008_));
 sky130_fd_sc_hd__xnor2_1 _15555_ (.A(_13085_),
    .B(_05008_),
    .Y(_05009_));
 sky130_fd_sc_hd__nand2_1 _15556_ (.A(\w[62][25] ),
    .B(net353),
    .Y(_05010_));
 sky130_fd_sc_hd__o21a_4 _15557_ (.A1(net353),
    .A2(_05009_),
    .B1(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1359 ();
 sky130_fd_sc_hd__nand2_1 _15559_ (.A(net746),
    .B(_04786_),
    .Y(_05013_));
 sky130_fd_sc_hd__o21ai_0 _15560_ (.A1(_04786_),
    .A2(_05011_),
    .B1(_05013_),
    .Y(_00146_));
 sky130_fd_sc_hd__nor3_1 _15561_ (.A(_13076_),
    .B(_13080_),
    .C(_13084_),
    .Y(_05014_));
 sky130_fd_sc_hd__or2_0 _15562_ (.A(_13081_),
    .B(_13080_),
    .X(_05015_));
 sky130_fd_sc_hd__a21oi_2 _15563_ (.A1(_13085_),
    .A2(_05015_),
    .B1(_13084_),
    .Y(_05016_));
 sky130_fd_sc_hd__a31oi_4 _15564_ (.A1(_04994_),
    .A2(_04996_),
    .A3(_05014_),
    .B1(_05016_),
    .Y(_05017_));
 sky130_fd_sc_hd__xnor2_2 _15565_ (.A(_13089_),
    .B(_05017_),
    .Y(_05018_));
 sky130_fd_sc_hd__nor2_1 _15566_ (.A(net353),
    .B(_05018_),
    .Y(_05019_));
 sky130_fd_sc_hd__a21oi_4 _15567_ (.A1(\w[62][26] ),
    .A2(net353),
    .B1(_05019_),
    .Y(_05020_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1358 ();
 sky130_fd_sc_hd__nand2_1 _15569_ (.A(net735),
    .B(_04786_),
    .Y(_05022_));
 sky130_fd_sc_hd__o21ai_0 _15570_ (.A1(_04786_),
    .A2(_05020_),
    .B1(_05022_),
    .Y(_00147_));
 sky130_fd_sc_hd__nand2_1 _15571_ (.A(_13085_),
    .B(_13089_),
    .Y(_05023_));
 sky130_fd_sc_hd__inv_1 _15572_ (.A(_13085_),
    .Y(_05024_));
 sky130_fd_sc_hd__o21bai_1 _15573_ (.A1(_05024_),
    .A2(_05007_),
    .B1_N(_13084_),
    .Y(_05025_));
 sky130_fd_sc_hd__a21oi_1 _15574_ (.A1(_13089_),
    .A2(_05025_),
    .B1(_13088_),
    .Y(_05026_));
 sky130_fd_sc_hd__o21ai_2 _15575_ (.A1(_05006_),
    .A2(_05023_),
    .B1(_05026_),
    .Y(_05027_));
 sky130_fd_sc_hd__xor2_4 _15576_ (.A(_13093_),
    .B(_05027_),
    .X(_05028_));
 sky130_fd_sc_hd__mux2i_4 _15577_ (.A0(\w[62][27] ),
    .A1(_05028_),
    .S(_04797_),
    .Y(_05029_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1357 ();
 sky130_fd_sc_hd__nand2_1 _15579_ (.A(net712),
    .B(_04786_),
    .Y(_05031_));
 sky130_fd_sc_hd__o21ai_0 _15580_ (.A1(_04786_),
    .A2(_05029_),
    .B1(_05031_),
    .Y(_00148_));
 sky130_fd_sc_hd__a21o_1 _15581_ (.A1(_13093_),
    .A2(_13088_),
    .B1(_13092_),
    .X(_05032_));
 sky130_fd_sc_hd__a31oi_2 _15582_ (.A1(_13089_),
    .A2(_13093_),
    .A3(_05017_),
    .B1(_05032_),
    .Y(_05033_));
 sky130_fd_sc_hd__xnor2_4 _15583_ (.A(_13097_),
    .B(_05033_),
    .Y(_05034_));
 sky130_fd_sc_hd__mux2i_4 _15584_ (.A0(\w[62][28] ),
    .A1(_05034_),
    .S(_04797_),
    .Y(_05035_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1356 ();
 sky130_fd_sc_hd__nand2_1 _15586_ (.A(net601),
    .B(_04786_),
    .Y(_05037_));
 sky130_fd_sc_hd__o21ai_0 _15587_ (.A1(_04786_),
    .A2(_05035_),
    .B1(_05037_),
    .Y(_00149_));
 sky130_fd_sc_hd__nand4_1 _15588_ (.A(_13085_),
    .B(_13089_),
    .C(_13093_),
    .D(_13097_),
    .Y(_05038_));
 sky130_fd_sc_hd__nor2b_1 _15589_ (.A(_05026_),
    .B_N(_13093_),
    .Y(_05039_));
 sky130_fd_sc_hd__o21a_1 _15590_ (.A1(_13092_),
    .A2(_05039_),
    .B1(_13097_),
    .X(_05040_));
 sky130_fd_sc_hd__nor2_2 _15591_ (.A(_13096_),
    .B(_05040_),
    .Y(_05041_));
 sky130_fd_sc_hd__o21ai_4 _15592_ (.A1(_05006_),
    .A2(_05038_),
    .B1(_05041_),
    .Y(_05042_));
 sky130_fd_sc_hd__xor2_4 _15593_ (.A(_13101_),
    .B(_05042_),
    .X(_05043_));
 sky130_fd_sc_hd__mux2i_4 _15594_ (.A0(\w[62][29] ),
    .A1(_05043_),
    .S(_04797_),
    .Y(_05044_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1355 ();
 sky130_fd_sc_hd__nand2_1 _15596_ (.A(net223),
    .B(_04786_),
    .Y(_05046_));
 sky130_fd_sc_hd__o21ai_0 _15597_ (.A1(_04786_),
    .A2(_05044_),
    .B1(_05046_),
    .Y(_00150_));
 sky130_fd_sc_hd__a21oi_2 _15598_ (.A1(_13089_),
    .A2(_05017_),
    .B1(_13088_),
    .Y(_05047_));
 sky130_fd_sc_hd__nand2_1 _15599_ (.A(_13097_),
    .B(_13101_),
    .Y(_05048_));
 sky130_fd_sc_hd__nor3_1 _15600_ (.A(_13105_),
    .B(net354),
    .C(_05048_),
    .Y(_05049_));
 sky130_fd_sc_hd__nand2_1 _15601_ (.A(_13093_),
    .B(_05049_),
    .Y(_05050_));
 sky130_fd_sc_hd__nand2b_1 _15602_ (.A_N(_13100_),
    .B(_13105_),
    .Y(_05051_));
 sky130_fd_sc_hd__nor3_1 _15603_ (.A(_13096_),
    .B(net354),
    .C(_05051_),
    .Y(_05052_));
 sky130_fd_sc_hd__nand3b_1 _15604_ (.A_N(_13092_),
    .B(_05047_),
    .C(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hd__o21ai_0 _15605_ (.A1(_13093_),
    .A2(_13092_),
    .B1(_13097_),
    .Y(_05054_));
 sky130_fd_sc_hd__a21oi_1 _15606_ (.A1(_13101_),
    .A2(_13096_),
    .B1(_13100_),
    .Y(_05055_));
 sky130_fd_sc_hd__o22a_1 _15607_ (.A1(_13105_),
    .A2(_05055_),
    .B1(_05051_),
    .B2(_13101_),
    .X(_05056_));
 sky130_fd_sc_hd__nand2_1 _15608_ (.A(\w[62][30] ),
    .B(net356),
    .Y(_05057_));
 sky130_fd_sc_hd__o21ai_0 _15609_ (.A1(net356),
    .A2(_05056_),
    .B1(_05057_),
    .Y(_05058_));
 sky130_fd_sc_hd__a221oi_1 _15610_ (.A1(_05052_),
    .A2(_05054_),
    .B1(_05049_),
    .B2(_13092_),
    .C1(_05058_),
    .Y(_05059_));
 sky130_fd_sc_hd__o211a_4 _15611_ (.A1(_05047_),
    .A2(_05050_),
    .B1(_05053_),
    .C1(_05059_),
    .X(_05060_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1354 ();
 sky130_fd_sc_hd__nand2_1 _15613_ (.A(net112),
    .B(_04786_),
    .Y(_05062_));
 sky130_fd_sc_hd__o21ai_0 _15614_ (.A1(_04786_),
    .A2(_05060_),
    .B1(_05062_),
    .Y(_00152_));
 sky130_fd_sc_hd__xor2_1 _15615_ (.A(_11822_),
    .B(_11825_),
    .X(_05063_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1350 ();
 sky130_fd_sc_hd__mux4_2 _15620_ (.A0(\w[0][31] ),
    .A1(\w[4][31] ),
    .A2(\w[2][31] ),
    .A3(\w[6][31] ),
    .S0(net481),
    .S1(net487),
    .X(_05068_));
 sky130_fd_sc_hd__mux4_2 _15621_ (.A0(\w[8][31] ),
    .A1(\w[12][31] ),
    .A2(\w[10][31] ),
    .A3(\w[14][31] ),
    .S0(net481),
    .S1(net487),
    .X(_05069_));
 sky130_fd_sc_hd__mux4_2 _15622_ (.A0(\w[16][31] ),
    .A1(\w[20][31] ),
    .A2(\w[18][31] ),
    .A3(\w[22][31] ),
    .S0(net481),
    .S1(net488),
    .X(_05070_));
 sky130_fd_sc_hd__mux4_2 _15623_ (.A0(\w[24][31] ),
    .A1(\w[28][31] ),
    .A2(\w[26][31] ),
    .A3(\w[30][31] ),
    .S0(net481),
    .S1(net488),
    .X(_05071_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1349 ();
 sky130_fd_sc_hd__mux4_2 _15625_ (.A0(_05068_),
    .A1(_05069_),
    .A2(_05070_),
    .A3(_05071_),
    .S0(net476),
    .S1(net475),
    .X(_05073_));
 sky130_fd_sc_hd__mux4_2 _15626_ (.A0(\w[32][31] ),
    .A1(\w[36][31] ),
    .A2(\w[34][31] ),
    .A3(\w[38][31] ),
    .S0(net481),
    .S1(net489),
    .X(_05074_));
 sky130_fd_sc_hd__mux4_2 _15627_ (.A0(\w[40][31] ),
    .A1(\w[44][31] ),
    .A2(\w[42][31] ),
    .A3(\w[46][31] ),
    .S0(net481),
    .S1(net489),
    .X(_05075_));
 sky130_fd_sc_hd__mux4_2 _15628_ (.A0(\w[48][31] ),
    .A1(\w[52][31] ),
    .A2(\w[50][31] ),
    .A3(\w[54][31] ),
    .S0(net481),
    .S1(net489),
    .X(_05076_));
 sky130_fd_sc_hd__mux4_2 _15629_ (.A0(\w[56][31] ),
    .A1(\w[60][31] ),
    .A2(\w[58][31] ),
    .A3(\w[62][31] ),
    .S0(net481),
    .S1(net489),
    .X(_05077_));
 sky130_fd_sc_hd__mux4_2 _15630_ (.A0(_05074_),
    .A1(_05075_),
    .A2(_05076_),
    .A3(_05077_),
    .S0(net476),
    .S1(net475),
    .X(_05078_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1348 ();
 sky130_fd_sc_hd__mux2i_4 _15632_ (.A0(_05073_),
    .A1(_05078_),
    .S(net473),
    .Y(_05080_));
 sky130_fd_sc_hd__xnor2_1 _15633_ (.A(_05063_),
    .B(_05080_),
    .Y(_05081_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1344 ();
 sky130_fd_sc_hd__mux4_2 _15638_ (.A0(\w[1][31] ),
    .A1(\w[5][31] ),
    .A2(\w[3][31] ),
    .A3(\w[7][31] ),
    .S0(net401),
    .S1(net409),
    .X(_05086_));
 sky130_fd_sc_hd__mux4_2 _15639_ (.A0(\w[9][31] ),
    .A1(\w[13][31] ),
    .A2(\w[11][31] ),
    .A3(\w[15][31] ),
    .S0(net401),
    .S1(net409),
    .X(_05087_));
 sky130_fd_sc_hd__mux4_2 _15640_ (.A0(\w[17][31] ),
    .A1(\w[21][31] ),
    .A2(\w[19][31] ),
    .A3(\w[23][31] ),
    .S0(net401),
    .S1(net409),
    .X(_05088_));
 sky130_fd_sc_hd__mux4_2 _15641_ (.A0(\w[25][31] ),
    .A1(\w[29][31] ),
    .A2(\w[27][31] ),
    .A3(\w[31][31] ),
    .S0(net401),
    .S1(net409),
    .X(_05089_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1343 ();
 sky130_fd_sc_hd__mux4_2 _15643_ (.A0(_05086_),
    .A1(_05087_),
    .A2(_05088_),
    .A3(_05089_),
    .S0(net400),
    .S1(net396),
    .X(_05091_));
 sky130_fd_sc_hd__mux4_2 _15644_ (.A0(\w[33][31] ),
    .A1(\w[37][31] ),
    .A2(\w[35][31] ),
    .A3(\w[39][31] ),
    .S0(net405),
    .S1(net409),
    .X(_05092_));
 sky130_fd_sc_hd__mux4_2 _15645_ (.A0(\w[41][31] ),
    .A1(\w[45][31] ),
    .A2(\w[43][31] ),
    .A3(\w[47][31] ),
    .S0(net405),
    .S1(net409),
    .X(_05093_));
 sky130_fd_sc_hd__mux4_2 _15646_ (.A0(\w[49][31] ),
    .A1(\w[53][31] ),
    .A2(\w[51][31] ),
    .A3(\w[55][31] ),
    .S0(net405),
    .S1(net409),
    .X(_05094_));
 sky130_fd_sc_hd__mux4_2 _15647_ (.A0(\w[57][31] ),
    .A1(\w[61][31] ),
    .A2(\w[59][31] ),
    .A3(\w[63][31] ),
    .S0(net405),
    .S1(net408),
    .X(_05095_));
 sky130_fd_sc_hd__mux4_2 _15648_ (.A0(_05092_),
    .A1(_05093_),
    .A2(_05094_),
    .A3(_05095_),
    .S0(net400),
    .S1(net536),
    .X(_05096_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1342 ();
 sky130_fd_sc_hd__mux2i_4 _15650_ (.A0(_05091_),
    .A1(_05096_),
    .S(net395),
    .Y(_05098_));
 sky130_fd_sc_hd__xnor2_4 _15651_ (.A(_11428_),
    .B(_05098_),
    .Y(_05099_));
 sky130_fd_sc_hd__xnor2_1 _15652_ (.A(_05081_),
    .B(_05099_),
    .Y(_05100_));
 sky130_fd_sc_hd__xor2_1 _15653_ (.A(_11104_),
    .B(_11300_),
    .X(_05101_));
 sky130_fd_sc_hd__xnor2_1 _15654_ (.A(_11006_),
    .B(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__xnor2_1 _15655_ (.A(_05100_),
    .B(_05102_),
    .Y(_05103_));
 sky130_fd_sc_hd__and2_4 _15656_ (.A(_04797_),
    .B(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__inv_1 _15657_ (.A(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__or3_4 _15658_ (.A(_13096_),
    .B(_13100_),
    .C(_05040_),
    .X(_05106_));
 sky130_fd_sc_hd__nor3_1 _15659_ (.A(_05004_),
    .B(_05005_),
    .C(_05106_),
    .Y(_05107_));
 sky130_fd_sc_hd__inv_1 _15660_ (.A(_05038_),
    .Y(_05108_));
 sky130_fd_sc_hd__o221ai_2 _15661_ (.A1(_13101_),
    .A2(_13100_),
    .B1(_05108_),
    .B2(_05106_),
    .C1(_13105_),
    .Y(_05109_));
 sky130_fd_sc_hd__nor3_1 _15662_ (.A(_13104_),
    .B(net354),
    .C(_05103_),
    .Y(_05110_));
 sky130_fd_sc_hd__o21ai_0 _15663_ (.A1(_05107_),
    .A2(_05109_),
    .B1(_05110_),
    .Y(_05111_));
 sky130_fd_sc_hd__o31a_1 _15664_ (.A1(_05105_),
    .A2(_05107_),
    .A3(_05109_),
    .B1(_05111_),
    .X(_05112_));
 sky130_fd_sc_hd__a22o_4 _15665_ (.A1(\w[62][31] ),
    .A2(net354),
    .B1(_05104_),
    .B2(_13104_),
    .X(_05113_));
 sky130_fd_sc_hd__mux2i_1 _15666_ (.A0(_05113_),
    .A1(net1),
    .S(_04786_),
    .Y(_05114_));
 sky130_fd_sc_hd__o21ai_0 _15667_ (.A1(_04786_),
    .A2(_05112_),
    .B1(_05114_),
    .Y(_00153_));
 sky130_fd_sc_hd__nor2b_4 _15668_ (.A(net1039),
    .B_N(_13536_),
    .Y(_05115_));
 sky130_fd_sc_hd__nand2_8 _15669_ (.A(_09797_),
    .B(_05115_),
    .Y(_05116_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1341 ();
 sky130_fd_sc_hd__mux2i_4 _15671_ (.A0(_13109_),
    .A1(\w[63][0] ),
    .S(net351),
    .Y(_05118_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1339 ();
 sky130_fd_sc_hd__nand2_1 _15674_ (.A(net739),
    .B(_05116_),
    .Y(_05121_));
 sky130_fd_sc_hd__o21ai_0 _15675_ (.A1(_05116_),
    .A2(_05118_),
    .B1(_05121_),
    .Y(_00353_));
 sky130_fd_sc_hd__mux2i_4 _15676_ (.A0(_13112_),
    .A1(\w[63][1] ),
    .S(net351),
    .Y(_05122_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1338 ();
 sky130_fd_sc_hd__nand2_1 _15678_ (.A(net738),
    .B(_05116_),
    .Y(_05124_));
 sky130_fd_sc_hd__o21ai_0 _15679_ (.A1(_05116_),
    .A2(_05122_),
    .B1(_05124_),
    .Y(_00364_));
 sky130_fd_sc_hd__nand2_4 _15680_ (.A(_11850_),
    .B(net339),
    .Y(_05125_));
 sky130_fd_sc_hd__o21ai_4 _15681_ (.A1(\w[63][2] ),
    .A2(net339),
    .B1(_05125_),
    .Y(_05126_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1337 ();
 sky130_fd_sc_hd__nand2_1 _15683_ (.A(net737),
    .B(_05116_),
    .Y(_05128_));
 sky130_fd_sc_hd__o21ai_0 _15684_ (.A1(_05116_),
    .A2(_05126_),
    .B1(_05128_),
    .Y(_00375_));
 sky130_fd_sc_hd__nor2b_2 _15685_ (.A(_13120_),
    .B_N(_11849_),
    .Y(_05129_));
 sky130_fd_sc_hd__nor2b_4 _15686_ (.A(_11849_),
    .B_N(_13120_),
    .Y(_05130_));
 sky130_fd_sc_hd__o21ai_4 _15687_ (.A1(_05129_),
    .A2(_05130_),
    .B1(net339),
    .Y(_05131_));
 sky130_fd_sc_hd__o21ai_4 _15688_ (.A1(\w[63][3] ),
    .A2(net339),
    .B1(_05131_),
    .Y(_05132_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1336 ();
 sky130_fd_sc_hd__nand2_1 _15690_ (.A(net736),
    .B(_05116_),
    .Y(_05134_));
 sky130_fd_sc_hd__o21ai_0 _15691_ (.A1(_05116_),
    .A2(_05132_),
    .B1(_05134_),
    .Y(_00378_));
 sky130_fd_sc_hd__inv_1 _15692_ (.A(_13124_),
    .Y(_05135_));
 sky130_fd_sc_hd__a21o_1 _15693_ (.A1(_13111_),
    .A2(_13116_),
    .B1(_13115_),
    .X(_05136_));
 sky130_fd_sc_hd__a21oi_1 _15694_ (.A1(_13120_),
    .A2(_05136_),
    .B1(_13119_),
    .Y(_05137_));
 sky130_fd_sc_hd__xnor2_1 _15695_ (.A(_05135_),
    .B(_05137_),
    .Y(_05138_));
 sky130_fd_sc_hd__nand2_2 _15696_ (.A(net339),
    .B(_05138_),
    .Y(_05139_));
 sky130_fd_sc_hd__o21ai_4 _15697_ (.A1(\w[63][4] ),
    .A2(net339),
    .B1(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1335 ();
 sky130_fd_sc_hd__nand2_1 _15699_ (.A(net734),
    .B(_05116_),
    .Y(_05142_));
 sky130_fd_sc_hd__o21ai_0 _15700_ (.A1(_05116_),
    .A2(_05140_),
    .B1(_05142_),
    .Y(_00379_));
 sky130_fd_sc_hd__inv_2 _15701_ (.A(_13123_),
    .Y(_05143_));
 sky130_fd_sc_hd__o21ai_2 _15702_ (.A1(_13119_),
    .A2(_05130_),
    .B1(_13124_),
    .Y(_05144_));
 sky130_fd_sc_hd__a21boi_4 _15703_ (.A1(_05143_),
    .A2(_05144_),
    .B1_N(_13128_),
    .Y(_05145_));
 sky130_fd_sc_hd__nand2_1 _15704_ (.A(_05143_),
    .B(_05144_),
    .Y(_05146_));
 sky130_fd_sc_hd__nor2_1 _15705_ (.A(_13128_),
    .B(_05146_),
    .Y(_05147_));
 sky130_fd_sc_hd__o21ai_4 _15706_ (.A1(_05145_),
    .A2(_05147_),
    .B1(net339),
    .Y(_05148_));
 sky130_fd_sc_hd__o21ai_4 _15707_ (.A1(\w[63][5] ),
    .A2(net339),
    .B1(_05148_),
    .Y(_05149_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1334 ();
 sky130_fd_sc_hd__nand2_1 _15709_ (.A(net733),
    .B(_05116_),
    .Y(_05151_));
 sky130_fd_sc_hd__o21ai_0 _15710_ (.A1(_05116_),
    .A2(_05149_),
    .B1(_05151_),
    .Y(_00380_));
 sky130_fd_sc_hd__inv_2 _15711_ (.A(_13132_),
    .Y(_05152_));
 sky130_fd_sc_hd__o21ai_1 _15712_ (.A1(_05135_),
    .A2(_05137_),
    .B1(_05143_),
    .Y(_05153_));
 sky130_fd_sc_hd__a21oi_2 _15713_ (.A1(_13128_),
    .A2(_05153_),
    .B1(_13127_),
    .Y(_05154_));
 sky130_fd_sc_hd__xnor2_1 _15714_ (.A(_05152_),
    .B(_05154_),
    .Y(_05155_));
 sky130_fd_sc_hd__nand2_2 _15715_ (.A(net339),
    .B(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__o21ai_4 _15716_ (.A1(\w[63][6] ),
    .A2(net339),
    .B1(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1333 ();
 sky130_fd_sc_hd__nand2_1 _15718_ (.A(net732),
    .B(_05116_),
    .Y(_05159_));
 sky130_fd_sc_hd__o21ai_0 _15719_ (.A1(_05116_),
    .A2(_05157_),
    .B1(_05159_),
    .Y(_00381_));
 sky130_fd_sc_hd__clkinv_2 _15720_ (.A(_13131_),
    .Y(_05160_));
 sky130_fd_sc_hd__o21ai_2 _15721_ (.A1(_13127_),
    .A2(_05145_),
    .B1(_13132_),
    .Y(_05161_));
 sky130_fd_sc_hd__a21boi_4 _15722_ (.A1(_05160_),
    .A2(_05161_),
    .B1_N(_13136_),
    .Y(_05162_));
 sky130_fd_sc_hd__nand2_1 _15723_ (.A(_05160_),
    .B(_05161_),
    .Y(_05163_));
 sky130_fd_sc_hd__nor2_1 _15724_ (.A(_13136_),
    .B(_05163_),
    .Y(_05164_));
 sky130_fd_sc_hd__o21ai_4 _15725_ (.A1(_05162_),
    .A2(_05164_),
    .B1(net339),
    .Y(_05165_));
 sky130_fd_sc_hd__o21ai_4 _15726_ (.A1(\w[63][7] ),
    .A2(net339),
    .B1(_05165_),
    .Y(_05166_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1332 ();
 sky130_fd_sc_hd__nand2_1 _15728_ (.A(net731),
    .B(_05116_),
    .Y(_05168_));
 sky130_fd_sc_hd__o21ai_0 _15729_ (.A1(_05116_),
    .A2(_05166_),
    .B1(_05168_),
    .Y(_00382_));
 sky130_fd_sc_hd__o21ai_2 _15730_ (.A1(_05152_),
    .A2(_05154_),
    .B1(_05160_),
    .Y(_05169_));
 sky130_fd_sc_hd__a21oi_1 _15731_ (.A1(_13136_),
    .A2(_05169_),
    .B1(_13135_),
    .Y(_05170_));
 sky130_fd_sc_hd__xor2_2 _15732_ (.A(_13140_),
    .B(_05170_),
    .X(_05171_));
 sky130_fd_sc_hd__nor2_1 _15733_ (.A(net350),
    .B(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__a21oi_4 _15734_ (.A1(\w[63][8] ),
    .A2(net350),
    .B1(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1331 ();
 sky130_fd_sc_hd__nand2_1 _15736_ (.A(net730),
    .B(_05116_),
    .Y(_05175_));
 sky130_fd_sc_hd__o21ai_0 _15737_ (.A1(_05116_),
    .A2(_05173_),
    .B1(_05175_),
    .Y(_00383_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1330 ();
 sky130_fd_sc_hd__inv_2 _15739_ (.A(_13139_),
    .Y(_05177_));
 sky130_fd_sc_hd__o21ai_2 _15740_ (.A1(_13135_),
    .A2(_05162_),
    .B1(_13140_),
    .Y(_05178_));
 sky130_fd_sc_hd__nand2_1 _15741_ (.A(_05177_),
    .B(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__and2_4 _15742_ (.A(_13144_),
    .B(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__nor2_1 _15743_ (.A(_13144_),
    .B(_05179_),
    .Y(_05181_));
 sky130_fd_sc_hd__o21ai_4 _15744_ (.A1(_05180_),
    .A2(_05181_),
    .B1(net339),
    .Y(_05182_));
 sky130_fd_sc_hd__o21ai_4 _15745_ (.A1(\w[63][9] ),
    .A2(net339),
    .B1(_05182_),
    .Y(_05183_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1329 ();
 sky130_fd_sc_hd__nand2_1 _15747_ (.A(net729),
    .B(_05116_),
    .Y(_05185_));
 sky130_fd_sc_hd__o21ai_0 _15748_ (.A1(_05116_),
    .A2(_05183_),
    .B1(_05185_),
    .Y(_00384_));
 sky130_fd_sc_hd__a211o_4 _15749_ (.A1(_13136_),
    .A2(_05169_),
    .B1(_13139_),
    .C1(_13135_),
    .X(_05186_));
 sky130_fd_sc_hd__o21ai_0 _15750_ (.A1(_13140_),
    .A2(_13139_),
    .B1(_13144_),
    .Y(_05187_));
 sky130_fd_sc_hd__inv_1 _15751_ (.A(_05187_),
    .Y(_05188_));
 sky130_fd_sc_hd__a21o_1 _15752_ (.A1(_05186_),
    .A2(_05188_),
    .B1(_13143_),
    .X(_05189_));
 sky130_fd_sc_hd__xnor2_1 _15753_ (.A(_13148_),
    .B(_05189_),
    .Y(_05190_));
 sky130_fd_sc_hd__nor2_4 _15754_ (.A(net355),
    .B(_05190_),
    .Y(_05191_));
 sky130_fd_sc_hd__a21oi_4 _15755_ (.A1(\w[63][10] ),
    .A2(net350),
    .B1(_05191_),
    .Y(_05192_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1327 ();
 sky130_fd_sc_hd__nand2_1 _15758_ (.A(net728),
    .B(_05116_),
    .Y(_05195_));
 sky130_fd_sc_hd__o21ai_0 _15759_ (.A1(_05116_),
    .A2(_05192_),
    .B1(_05195_),
    .Y(_00354_));
 sky130_fd_sc_hd__nand3_2 _15760_ (.A(_13144_),
    .B(_13148_),
    .C(_13152_),
    .Y(_05196_));
 sky130_fd_sc_hd__a21oi_4 _15761_ (.A1(_05177_),
    .A2(_05178_),
    .B1(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__a21oi_1 _15762_ (.A1(_13148_),
    .A2(_13143_),
    .B1(_13147_),
    .Y(_05198_));
 sky130_fd_sc_hd__nor2b_4 _15763_ (.A(_05198_),
    .B_N(_13152_),
    .Y(_05199_));
 sky130_fd_sc_hd__nor2_4 _15764_ (.A(_05197_),
    .B(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__o21ai_0 _15765_ (.A1(_13143_),
    .A2(_05180_),
    .B1(_13148_),
    .Y(_05201_));
 sky130_fd_sc_hd__or3b_1 _15766_ (.A(_13152_),
    .B(_13147_),
    .C_N(_05201_),
    .X(_05202_));
 sky130_fd_sc_hd__and3_4 _15767_ (.A(net339),
    .B(_05200_),
    .C(_05202_),
    .X(_05203_));
 sky130_fd_sc_hd__a21oi_4 _15768_ (.A1(\w[63][11] ),
    .A2(net352),
    .B1(_05203_),
    .Y(_05204_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1326 ();
 sky130_fd_sc_hd__nand2_1 _15770_ (.A(net727),
    .B(_05116_),
    .Y(_05206_));
 sky130_fd_sc_hd__o21ai_0 _15771_ (.A1(_05116_),
    .A2(_05204_),
    .B1(_05206_),
    .Y(_00355_));
 sky130_fd_sc_hd__inv_1 _15772_ (.A(_13156_),
    .Y(_05207_));
 sky130_fd_sc_hd__a2111oi_2 _15773_ (.A1(_05186_),
    .A2(_05188_),
    .B1(_13143_),
    .C1(_13147_),
    .D1(_13151_),
    .Y(_05208_));
 sky130_fd_sc_hd__or2_0 _15774_ (.A(_13148_),
    .B(_13147_),
    .X(_05209_));
 sky130_fd_sc_hd__a21oi_2 _15775_ (.A1(_13152_),
    .A2(_05209_),
    .B1(_13151_),
    .Y(_05210_));
 sky130_fd_sc_hd__or2_4 _15776_ (.A(_05208_),
    .B(_05210_),
    .X(_05211_));
 sky130_fd_sc_hd__xnor2_1 _15777_ (.A(_05207_),
    .B(_05211_),
    .Y(_05212_));
 sky130_fd_sc_hd__nand2_2 _15778_ (.A(net339),
    .B(_05212_),
    .Y(_05213_));
 sky130_fd_sc_hd__o21ai_4 _15779_ (.A1(\w[63][12] ),
    .A2(net339),
    .B1(_05213_),
    .Y(_05214_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1325 ();
 sky130_fd_sc_hd__nand2_1 _15781_ (.A(net726),
    .B(_05116_),
    .Y(_05216_));
 sky130_fd_sc_hd__o21ai_0 _15782_ (.A1(_05116_),
    .A2(_05214_),
    .B1(_05216_),
    .Y(_00356_));
 sky130_fd_sc_hd__or3_1 _15783_ (.A(_13151_),
    .B(_05197_),
    .C(_05199_),
    .X(_05217_));
 sky130_fd_sc_hd__a21oi_1 _15784_ (.A1(_13156_),
    .A2(_05217_),
    .B1(_13155_),
    .Y(_05218_));
 sky130_fd_sc_hd__xor2_1 _15785_ (.A(_13160_),
    .B(_05218_),
    .X(_05219_));
 sky130_fd_sc_hd__nor2_1 _15786_ (.A(net355),
    .B(_05219_),
    .Y(_05220_));
 sky130_fd_sc_hd__a21oi_4 _15787_ (.A1(\w[63][13] ),
    .A2(net355),
    .B1(_05220_),
    .Y(_05221_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1324 ();
 sky130_fd_sc_hd__nand2_1 _15789_ (.A(net723),
    .B(_05116_),
    .Y(_05223_));
 sky130_fd_sc_hd__o21ai_0 _15790_ (.A1(_05116_),
    .A2(_05221_),
    .B1(_05223_),
    .Y(_00357_));
 sky130_fd_sc_hd__o21bai_1 _15791_ (.A1(_05207_),
    .A2(_05211_),
    .B1_N(_13155_),
    .Y(_05224_));
 sky130_fd_sc_hd__a21oi_1 _15792_ (.A1(_13160_),
    .A2(_05224_),
    .B1(_13159_),
    .Y(_05225_));
 sky130_fd_sc_hd__xor2_2 _15793_ (.A(_13164_),
    .B(_05225_),
    .X(_05226_));
 sky130_fd_sc_hd__nor2_2 _15794_ (.A(net350),
    .B(_05226_),
    .Y(_05227_));
 sky130_fd_sc_hd__a21oi_4 _15795_ (.A1(\w[63][14] ),
    .A2(net350),
    .B1(_05227_),
    .Y(_05228_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1323 ();
 sky130_fd_sc_hd__nand2_1 _15797_ (.A(net711),
    .B(_05116_),
    .Y(_05230_));
 sky130_fd_sc_hd__o21ai_0 _15798_ (.A1(_05116_),
    .A2(_05228_),
    .B1(_05230_),
    .Y(_00358_));
 sky130_fd_sc_hd__nand3_2 _15799_ (.A(_13156_),
    .B(_13160_),
    .C(_13164_),
    .Y(_05231_));
 sky130_fd_sc_hd__a21o_1 _15800_ (.A1(_13156_),
    .A2(_13151_),
    .B1(_13155_),
    .X(_05232_));
 sky130_fd_sc_hd__a21o_1 _15801_ (.A1(_13160_),
    .A2(_05232_),
    .B1(_13159_),
    .X(_05233_));
 sky130_fd_sc_hd__a21oi_1 _15802_ (.A1(_13164_),
    .A2(_05233_),
    .B1(_13163_),
    .Y(_05234_));
 sky130_fd_sc_hd__o21ai_2 _15803_ (.A1(_05200_),
    .A2(_05231_),
    .B1(_05234_),
    .Y(_05235_));
 sky130_fd_sc_hd__xnor2_2 _15804_ (.A(_13168_),
    .B(_05235_),
    .Y(_05236_));
 sky130_fd_sc_hd__nand2_4 _15805_ (.A(net339),
    .B(_05236_),
    .Y(_05237_));
 sky130_fd_sc_hd__o21ai_4 _15806_ (.A1(\w[63][15] ),
    .A2(net339),
    .B1(_05237_),
    .Y(_05238_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1322 ();
 sky130_fd_sc_hd__nand2_1 _15808_ (.A(net700),
    .B(_05116_),
    .Y(_05240_));
 sky130_fd_sc_hd__o21ai_0 _15809_ (.A1(_05116_),
    .A2(_05238_),
    .B1(_05240_),
    .Y(_00359_));
 sky130_fd_sc_hd__a21o_1 _15810_ (.A1(_13160_),
    .A2(_13155_),
    .B1(_13159_),
    .X(_05241_));
 sky130_fd_sc_hd__a21oi_1 _15811_ (.A1(_13164_),
    .A2(_05241_),
    .B1(_13163_),
    .Y(_05242_));
 sky130_fd_sc_hd__o21ai_0 _15812_ (.A1(_05211_),
    .A2(_05231_),
    .B1(_05242_),
    .Y(_05243_));
 sky130_fd_sc_hd__a21oi_1 _15813_ (.A1(_13168_),
    .A2(_05243_),
    .B1(_13167_),
    .Y(_05244_));
 sky130_fd_sc_hd__xor2_1 _15814_ (.A(_13172_),
    .B(_05244_),
    .X(_05245_));
 sky130_fd_sc_hd__nor2_2 _15815_ (.A(net351),
    .B(_05245_),
    .Y(_05246_));
 sky130_fd_sc_hd__a21oi_4 _15816_ (.A1(\w[63][16] ),
    .A2(net351),
    .B1(_05246_),
    .Y(_05247_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1321 ();
 sky130_fd_sc_hd__nand2_1 _15818_ (.A(net689),
    .B(_05116_),
    .Y(_05249_));
 sky130_fd_sc_hd__o21ai_0 _15819_ (.A1(_05116_),
    .A2(_05247_),
    .B1(_05249_),
    .Y(_00360_));
 sky130_fd_sc_hd__nand2_1 _15820_ (.A(_13168_),
    .B(_13172_),
    .Y(_05250_));
 sky130_fd_sc_hd__or2_4 _15821_ (.A(_05231_),
    .B(_05250_),
    .X(_05251_));
 sky130_fd_sc_hd__inv_1 _15822_ (.A(_13168_),
    .Y(_05252_));
 sky130_fd_sc_hd__o21bai_1 _15823_ (.A1(_05252_),
    .A2(_05234_),
    .B1_N(_13167_),
    .Y(_05253_));
 sky130_fd_sc_hd__a21oi_2 _15824_ (.A1(_13172_),
    .A2(_05253_),
    .B1(_13171_),
    .Y(_05254_));
 sky130_fd_sc_hd__o21ai_2 _15825_ (.A1(_05200_),
    .A2(_05251_),
    .B1(_05254_),
    .Y(_05255_));
 sky130_fd_sc_hd__xnor2_4 _15826_ (.A(_13176_),
    .B(_05255_),
    .Y(_05256_));
 sky130_fd_sc_hd__nand2_2 _15827_ (.A(net339),
    .B(_05256_),
    .Y(_05257_));
 sky130_fd_sc_hd__o21ai_4 _15828_ (.A1(\w[63][17] ),
    .A2(net339),
    .B1(_05257_),
    .Y(_05258_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1320 ();
 sky130_fd_sc_hd__nand2_1 _15830_ (.A(net678),
    .B(_05116_),
    .Y(_05260_));
 sky130_fd_sc_hd__o21ai_0 _15831_ (.A1(_05116_),
    .A2(_05258_),
    .B1(_05260_),
    .Y(_00361_));
 sky130_fd_sc_hd__o21bai_1 _15832_ (.A1(_05252_),
    .A2(_05242_),
    .B1_N(_13167_),
    .Y(_05261_));
 sky130_fd_sc_hd__a21oi_2 _15833_ (.A1(_13172_),
    .A2(_05261_),
    .B1(_13171_),
    .Y(_05262_));
 sky130_fd_sc_hd__o21ai_0 _15834_ (.A1(_05211_),
    .A2(_05251_),
    .B1(_05262_),
    .Y(_05263_));
 sky130_fd_sc_hd__a21oi_1 _15835_ (.A1(_13176_),
    .A2(_05263_),
    .B1(_13175_),
    .Y(_05264_));
 sky130_fd_sc_hd__xor2_1 _15836_ (.A(_13180_),
    .B(_05264_),
    .X(_05265_));
 sky130_fd_sc_hd__nor2_2 _15837_ (.A(net350),
    .B(_05265_),
    .Y(_05266_));
 sky130_fd_sc_hd__a21oi_4 _15838_ (.A1(\w[63][18] ),
    .A2(net350),
    .B1(_05266_),
    .Y(_05267_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1319 ();
 sky130_fd_sc_hd__nand2_1 _15840_ (.A(net667),
    .B(_05116_),
    .Y(_05269_));
 sky130_fd_sc_hd__o21ai_0 _15841_ (.A1(_05116_),
    .A2(_05267_),
    .B1(_05269_),
    .Y(_00362_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1318 ();
 sky130_fd_sc_hd__nand2_2 _15843_ (.A(_13176_),
    .B(_13180_),
    .Y(_05271_));
 sky130_fd_sc_hd__nor2_2 _15844_ (.A(_05251_),
    .B(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__o21ai_4 _15845_ (.A1(_05197_),
    .A2(_05199_),
    .B1(_05272_),
    .Y(_05273_));
 sky130_fd_sc_hd__nor2_2 _15846_ (.A(_05254_),
    .B(_05271_),
    .Y(_05274_));
 sky130_fd_sc_hd__a21oi_4 _15847_ (.A1(_13180_),
    .A2(_13175_),
    .B1(_05274_),
    .Y(_05275_));
 sky130_fd_sc_hd__nand2_1 _15848_ (.A(_05273_),
    .B(_05275_),
    .Y(_05276_));
 sky130_fd_sc_hd__nor2_1 _15849_ (.A(_13179_),
    .B(_05276_),
    .Y(_05277_));
 sky130_fd_sc_hd__xor2_1 _15850_ (.A(_13184_),
    .B(_05277_),
    .X(_05278_));
 sky130_fd_sc_hd__nor2_1 _15851_ (.A(net355),
    .B(_05278_),
    .Y(_05279_));
 sky130_fd_sc_hd__a21oi_4 _15852_ (.A1(\w[63][19] ),
    .A2(net355),
    .B1(_05279_),
    .Y(_05280_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1317 ();
 sky130_fd_sc_hd__nand2_1 _15854_ (.A(net656),
    .B(_05116_),
    .Y(_05282_));
 sky130_fd_sc_hd__o21ai_0 _15855_ (.A1(_05116_),
    .A2(_05280_),
    .B1(_05282_),
    .Y(_00363_));
 sky130_fd_sc_hd__o21a_1 _15856_ (.A1(_13176_),
    .A2(_13175_),
    .B1(_13180_),
    .X(_05283_));
 sky130_fd_sc_hd__o21ai_2 _15857_ (.A1(_13179_),
    .A2(_05283_),
    .B1(_13184_),
    .Y(_05284_));
 sky130_fd_sc_hd__nand2b_4 _15858_ (.A_N(_13183_),
    .B(_05284_),
    .Y(_05285_));
 sky130_fd_sc_hd__nor3_1 _15859_ (.A(_13175_),
    .B(_13179_),
    .C(_13183_),
    .Y(_05286_));
 sky130_fd_sc_hd__o311ai_4 _15860_ (.A1(_05208_),
    .A2(_05210_),
    .A3(_05251_),
    .B1(_05262_),
    .C1(_05286_),
    .Y(_05287_));
 sky130_fd_sc_hd__and3_1 _15861_ (.A(_13188_),
    .B(_05285_),
    .C(_05287_),
    .X(_05288_));
 sky130_fd_sc_hd__a21oi_1 _15862_ (.A1(_05285_),
    .A2(_05287_),
    .B1(_13188_),
    .Y(_05289_));
 sky130_fd_sc_hd__o21ai_2 _15863_ (.A1(_05288_),
    .A2(_05289_),
    .B1(net339),
    .Y(_05290_));
 sky130_fd_sc_hd__o21ai_4 _15864_ (.A1(\w[63][20] ),
    .A2(net339),
    .B1(_05290_),
    .Y(_05291_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1315 ();
 sky130_fd_sc_hd__nand2_1 _15867_ (.A(net645),
    .B(_05116_),
    .Y(_05294_));
 sky130_fd_sc_hd__o21ai_0 _15868_ (.A1(_05116_),
    .A2(_05291_),
    .B1(_05294_),
    .Y(_00365_));
 sky130_fd_sc_hd__nor2_1 _15869_ (.A(_13179_),
    .B(_13183_),
    .Y(_05295_));
 sky130_fd_sc_hd__o21ai_0 _15870_ (.A1(_13184_),
    .A2(_13183_),
    .B1(_13188_),
    .Y(_05296_));
 sky130_fd_sc_hd__a31oi_1 _15871_ (.A1(_05273_),
    .A2(_05275_),
    .A3(_05295_),
    .B1(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__nor2_1 _15872_ (.A(_13187_),
    .B(_05297_),
    .Y(_05298_));
 sky130_fd_sc_hd__xor2_2 _15873_ (.A(_13192_),
    .B(_05298_),
    .X(_05299_));
 sky130_fd_sc_hd__nor2_2 _15874_ (.A(net350),
    .B(_05299_),
    .Y(_05300_));
 sky130_fd_sc_hd__a21oi_4 _15875_ (.A1(\w[63][21] ),
    .A2(net350),
    .B1(_05300_),
    .Y(_05301_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1314 ();
 sky130_fd_sc_hd__nand2_1 _15877_ (.A(net634),
    .B(_05116_),
    .Y(_05303_));
 sky130_fd_sc_hd__o21ai_0 _15878_ (.A1(_05116_),
    .A2(_05301_),
    .B1(_05303_),
    .Y(_00366_));
 sky130_fd_sc_hd__clkinv_1 _15879_ (.A(_13196_),
    .Y(_05304_));
 sky130_fd_sc_hd__a21o_4 _15880_ (.A1(_13192_),
    .A2(_13187_),
    .B1(_13191_),
    .X(_05305_));
 sky130_fd_sc_hd__a41oi_4 _15881_ (.A1(_13188_),
    .A2(_13192_),
    .A3(_05285_),
    .A4(_05287_),
    .B1(_05305_),
    .Y(_05306_));
 sky130_fd_sc_hd__xnor2_2 _15882_ (.A(_05304_),
    .B(_05306_),
    .Y(_05307_));
 sky130_fd_sc_hd__nand2_2 _15883_ (.A(net339),
    .B(_05307_),
    .Y(_05308_));
 sky130_fd_sc_hd__o21ai_4 _15884_ (.A1(\w[63][22] ),
    .A2(net339),
    .B1(_05308_),
    .Y(_05309_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1313 ();
 sky130_fd_sc_hd__nand2_1 _15886_ (.A(net623),
    .B(_05116_),
    .Y(_05311_));
 sky130_fd_sc_hd__o21ai_0 _15887_ (.A1(_05116_),
    .A2(_05309_),
    .B1(_05311_),
    .Y(_00367_));
 sky130_fd_sc_hd__nor3_2 _15888_ (.A(_13179_),
    .B(_13183_),
    .C(_05305_),
    .Y(_05312_));
 sky130_fd_sc_hd__nand2b_1 _15889_ (.A_N(_13187_),
    .B(_05296_),
    .Y(_05313_));
 sky130_fd_sc_hd__a21o_4 _15890_ (.A1(_13192_),
    .A2(_05313_),
    .B1(_13191_),
    .X(_05314_));
 sky130_fd_sc_hd__nand2_1 _15891_ (.A(_13196_),
    .B(_05314_),
    .Y(_05315_));
 sky130_fd_sc_hd__a31oi_2 _15892_ (.A1(_05273_),
    .A2(_05275_),
    .A3(_05312_),
    .B1(_05315_),
    .Y(_05316_));
 sky130_fd_sc_hd__o21a_4 _15893_ (.A1(_13195_),
    .A2(_05316_),
    .B1(_13200_),
    .X(_05317_));
 sky130_fd_sc_hd__nor3_1 _15894_ (.A(_13200_),
    .B(_13195_),
    .C(_05316_),
    .Y(_05318_));
 sky130_fd_sc_hd__o21ai_4 _15895_ (.A1(_05317_),
    .A2(_05318_),
    .B1(net339),
    .Y(_05319_));
 sky130_fd_sc_hd__o21ai_4 _15896_ (.A1(\w[63][23] ),
    .A2(net339),
    .B1(_05319_),
    .Y(_05320_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1312 ();
 sky130_fd_sc_hd__nand2_1 _15898_ (.A(net612),
    .B(_05116_),
    .Y(_05322_));
 sky130_fd_sc_hd__o21ai_0 _15899_ (.A1(_05116_),
    .A2(_05320_),
    .B1(_05322_),
    .Y(_00368_));
 sky130_fd_sc_hd__o21bai_1 _15900_ (.A1(_05304_),
    .A2(_05306_),
    .B1_N(_13195_),
    .Y(_05323_));
 sky130_fd_sc_hd__a21oi_2 _15901_ (.A1(_13200_),
    .A2(_05323_),
    .B1(_13199_),
    .Y(_05324_));
 sky130_fd_sc_hd__xnor2_2 _15902_ (.A(_13204_),
    .B(_05324_),
    .Y(_05325_));
 sky130_fd_sc_hd__mux2i_4 _15903_ (.A0(\w[63][24] ),
    .A1(_05325_),
    .S(net339),
    .Y(_05326_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1311 ();
 sky130_fd_sc_hd__nand2_1 _15905_ (.A(net600),
    .B(_05116_),
    .Y(_05328_));
 sky130_fd_sc_hd__o21ai_0 _15906_ (.A1(_05116_),
    .A2(net1145),
    .B1(_05328_),
    .Y(_00369_));
 sky130_fd_sc_hd__o21ai_2 _15907_ (.A1(_13199_),
    .A2(_05317_),
    .B1(_13204_),
    .Y(_05329_));
 sky130_fd_sc_hd__nor2_2 _15908_ (.A(_13208_),
    .B(_13203_),
    .Y(_05330_));
 sky130_fd_sc_hd__a21o_1 _15909_ (.A1(_13200_),
    .A2(_13195_),
    .B1(_13199_),
    .X(_05331_));
 sky130_fd_sc_hd__a21o_4 _15910_ (.A1(_13204_),
    .A2(_05331_),
    .B1(_13203_),
    .X(_05332_));
 sky130_fd_sc_hd__and3_4 _15911_ (.A(_13196_),
    .B(_13200_),
    .C(_13204_),
    .X(_05333_));
 sky130_fd_sc_hd__nand2_1 _15912_ (.A(_05314_),
    .B(_05333_),
    .Y(_05334_));
 sky130_fd_sc_hd__a31oi_1 _15913_ (.A1(_05273_),
    .A2(_05275_),
    .A3(_05312_),
    .B1(_05334_),
    .Y(_05335_));
 sky130_fd_sc_hd__o21ai_0 _15914_ (.A1(_05332_),
    .A2(_05335_),
    .B1(_13208_),
    .Y(_05336_));
 sky130_fd_sc_hd__nand2_2 _15915_ (.A(net339),
    .B(_05336_),
    .Y(_05337_));
 sky130_fd_sc_hd__a21oi_4 _15916_ (.A1(_05329_),
    .A2(_05330_),
    .B1(_05337_),
    .Y(_05338_));
 sky130_fd_sc_hd__a21oi_4 _15917_ (.A1(\w[63][25] ),
    .A2(net350),
    .B1(_05338_),
    .Y(_05339_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1310 ();
 sky130_fd_sc_hd__nand2_1 _15919_ (.A(net589),
    .B(_05116_),
    .Y(_05341_));
 sky130_fd_sc_hd__o21ai_0 _15920_ (.A1(_05116_),
    .A2(_05339_),
    .B1(_05341_),
    .Y(_00370_));
 sky130_fd_sc_hd__nand2_2 _15921_ (.A(_13208_),
    .B(_05333_),
    .Y(_05342_));
 sky130_fd_sc_hd__a21oi_1 _15922_ (.A1(_13208_),
    .A2(_05332_),
    .B1(_13207_),
    .Y(_05343_));
 sky130_fd_sc_hd__o21ai_2 _15923_ (.A1(_05306_),
    .A2(_05342_),
    .B1(_05343_),
    .Y(_05344_));
 sky130_fd_sc_hd__xnor2_1 _15924_ (.A(_13212_),
    .B(_05344_),
    .Y(_05345_));
 sky130_fd_sc_hd__nand2_2 _15925_ (.A(net339),
    .B(_05345_),
    .Y(_05346_));
 sky130_fd_sc_hd__o21ai_4 _15926_ (.A1(\w[63][26] ),
    .A2(net339),
    .B1(_05346_),
    .Y(_05347_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1309 ();
 sky130_fd_sc_hd__nand2_1 _15928_ (.A(net578),
    .B(_05116_),
    .Y(_05349_));
 sky130_fd_sc_hd__o21ai_0 _15929_ (.A1(_05116_),
    .A2(_05347_),
    .B1(_05349_),
    .Y(_00371_));
 sky130_fd_sc_hd__inv_1 _15930_ (.A(_13212_),
    .Y(_05350_));
 sky130_fd_sc_hd__nand3_2 _15931_ (.A(_05273_),
    .B(_05275_),
    .C(_05312_),
    .Y(_05351_));
 sky130_fd_sc_hd__nor2b_2 _15932_ (.A(_05342_),
    .B_N(_05314_),
    .Y(_05352_));
 sky130_fd_sc_hd__a21boi_4 _15933_ (.A1(_05351_),
    .A2(_05352_),
    .B1_N(_05343_),
    .Y(_05353_));
 sky130_fd_sc_hd__o21bai_1 _15934_ (.A1(_05350_),
    .A2(_05353_),
    .B1_N(_13211_),
    .Y(_05354_));
 sky130_fd_sc_hd__nor2_1 _15935_ (.A(_13216_),
    .B(_05354_),
    .Y(_05355_));
 sky130_fd_sc_hd__and2_0 _15936_ (.A(_13216_),
    .B(_05354_),
    .X(_05356_));
 sky130_fd_sc_hd__nand2_1 _15937_ (.A(\w[63][27] ),
    .B(net351),
    .Y(_05357_));
 sky130_fd_sc_hd__o31a_2 _15938_ (.A1(net351),
    .A2(_05355_),
    .A3(_05356_),
    .B1(_05357_),
    .X(_05358_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1308 ();
 sky130_fd_sc_hd__nand2_1 _15940_ (.A(net567),
    .B(_05116_),
    .Y(_05360_));
 sky130_fd_sc_hd__o21ai_0 _15941_ (.A1(_05116_),
    .A2(_05358_),
    .B1(_05360_),
    .Y(_00372_));
 sky130_fd_sc_hd__and4_4 _15942_ (.A(_13188_),
    .B(_13192_),
    .C(_13208_),
    .D(_05333_),
    .X(_05361_));
 sky130_fd_sc_hd__nand2_1 _15943_ (.A(_13208_),
    .B(_05332_),
    .Y(_05362_));
 sky130_fd_sc_hd__nand3_1 _15944_ (.A(_13208_),
    .B(_05305_),
    .C(_05333_),
    .Y(_05363_));
 sky130_fd_sc_hd__nand2_2 _15945_ (.A(_05362_),
    .B(_05363_),
    .Y(_05364_));
 sky130_fd_sc_hd__or3_4 _15946_ (.A(_13207_),
    .B(_13211_),
    .C(_13215_),
    .X(_05365_));
 sky130_fd_sc_hd__a311oi_4 _15947_ (.A1(_05285_),
    .A2(_05287_),
    .A3(_05361_),
    .B1(_05364_),
    .C1(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__or2_0 _15948_ (.A(_13212_),
    .B(_13211_),
    .X(_05367_));
 sky130_fd_sc_hd__a21oi_1 _15949_ (.A1(_13216_),
    .A2(_05367_),
    .B1(_13215_),
    .Y(_05368_));
 sky130_fd_sc_hd__nor2_1 _15950_ (.A(_05366_),
    .B(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__xnor2_1 _15951_ (.A(_13220_),
    .B(_05369_),
    .Y(_05370_));
 sky130_fd_sc_hd__nor2_4 _15952_ (.A(net351),
    .B(_05370_),
    .Y(_05371_));
 sky130_fd_sc_hd__a21oi_4 _15953_ (.A1(\w[63][28] ),
    .A2(done),
    .B1(_05371_),
    .Y(_05372_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1307 ();
 sky130_fd_sc_hd__nand2_1 _15955_ (.A(net556),
    .B(_05116_),
    .Y(_05374_));
 sky130_fd_sc_hd__o21ai_0 _15956_ (.A1(_05116_),
    .A2(_05372_),
    .B1(_05374_),
    .Y(_00373_));
 sky130_fd_sc_hd__nand3_1 _15957_ (.A(_13212_),
    .B(_13216_),
    .C(_13220_),
    .Y(_05375_));
 sky130_fd_sc_hd__a21o_1 _15958_ (.A1(_13216_),
    .A2(_13211_),
    .B1(_13215_),
    .X(_05376_));
 sky130_fd_sc_hd__a21oi_1 _15959_ (.A1(_13220_),
    .A2(_05376_),
    .B1(_13219_),
    .Y(_05377_));
 sky130_fd_sc_hd__o21ai_0 _15960_ (.A1(_05353_),
    .A2(_05375_),
    .B1(_05377_),
    .Y(_05378_));
 sky130_fd_sc_hd__xor2_1 _15961_ (.A(_13224_),
    .B(_05378_),
    .X(_05379_));
 sky130_fd_sc_hd__mux2i_4 _15962_ (.A0(\w[63][29] ),
    .A1(_05379_),
    .S(net339),
    .Y(_05380_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1306 ();
 sky130_fd_sc_hd__nand2_1 _15964_ (.A(net278),
    .B(_05116_),
    .Y(_05382_));
 sky130_fd_sc_hd__o21ai_0 _15965_ (.A1(_05116_),
    .A2(_05380_),
    .B1(_05382_),
    .Y(_00374_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1305 ();
 sky130_fd_sc_hd__nand2_1 _15967_ (.A(_13220_),
    .B(_13224_),
    .Y(_05384_));
 sky130_fd_sc_hd__a21oi_1 _15968_ (.A1(_13224_),
    .A2(_13219_),
    .B1(_13223_),
    .Y(_05385_));
 sky130_fd_sc_hd__o31ai_1 _15969_ (.A1(_05366_),
    .A2(_05368_),
    .A3(_05384_),
    .B1(_05385_),
    .Y(_05386_));
 sky130_fd_sc_hd__xnor2_1 _15970_ (.A(_13228_),
    .B(_05386_),
    .Y(_05387_));
 sky130_fd_sc_hd__nor2_2 _15971_ (.A(net351),
    .B(_05387_),
    .Y(_05388_));
 sky130_fd_sc_hd__a21oi_4 _15972_ (.A1(\w[63][30] ),
    .A2(net355),
    .B1(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__a21oi_1 _15973_ (.A1(_09797_),
    .A2(_05115_),
    .B1(net267),
    .Y(_05390_));
 sky130_fd_sc_hd__a31oi_1 _15974_ (.A1(_09797_),
    .A2(_05115_),
    .A3(net1143),
    .B1(_05390_),
    .Y(_00376_));
 sky130_fd_sc_hd__nand2_1 _15975_ (.A(_13220_),
    .B(_05376_),
    .Y(_05391_));
 sky130_fd_sc_hd__nor3_1 _15976_ (.A(_13219_),
    .B(_13223_),
    .C(_13227_),
    .Y(_05392_));
 sky130_fd_sc_hd__o211ai_1 _15977_ (.A1(_05353_),
    .A2(_05375_),
    .B1(_05391_),
    .C1(_05392_),
    .Y(_05393_));
 sky130_fd_sc_hd__nor3_1 _15978_ (.A(_13224_),
    .B(_13223_),
    .C(_13227_),
    .Y(_05394_));
 sky130_fd_sc_hd__nor2_1 _15979_ (.A(_13228_),
    .B(_13227_),
    .Y(_05395_));
 sky130_fd_sc_hd__nor2_1 _15980_ (.A(_05394_),
    .B(_05395_),
    .Y(_05396_));
 sky130_fd_sc_hd__xor2_1 _15981_ (.A(_12070_),
    .B(_12073_),
    .X(_05397_));
 sky130_fd_sc_hd__mux4_2 _15982_ (.A0(\w[1][31] ),
    .A1(\w[5][31] ),
    .A2(\w[3][31] ),
    .A3(\w[7][31] ),
    .S0(net459),
    .S1(net544),
    .X(_05398_));
 sky130_fd_sc_hd__mux4_2 _15983_ (.A0(\w[9][31] ),
    .A1(\w[13][31] ),
    .A2(\w[11][31] ),
    .A3(\w[15][31] ),
    .S0(net459),
    .S1(net544),
    .X(_05399_));
 sky130_fd_sc_hd__mux4_2 _15984_ (.A0(\w[17][31] ),
    .A1(\w[21][31] ),
    .A2(\w[19][31] ),
    .A3(\w[23][31] ),
    .S0(net459),
    .S1(net544),
    .X(_05400_));
 sky130_fd_sc_hd__mux4_2 _15985_ (.A0(\w[25][31] ),
    .A1(\w[29][31] ),
    .A2(\w[27][31] ),
    .A3(\w[31][31] ),
    .S0(net459),
    .S1(net544),
    .X(_05401_));
 sky130_fd_sc_hd__mux4_2 _15986_ (.A0(_05398_),
    .A1(_05399_),
    .A2(_05400_),
    .A3(_05401_),
    .S0(net456),
    .S1(net454),
    .X(_05402_));
 sky130_fd_sc_hd__mux4_2 _15987_ (.A0(\w[33][31] ),
    .A1(\w[37][31] ),
    .A2(\w[35][31] ),
    .A3(\w[39][31] ),
    .S0(net459),
    .S1(net470),
    .X(_05403_));
 sky130_fd_sc_hd__mux4_2 _15988_ (.A0(\w[41][31] ),
    .A1(\w[45][31] ),
    .A2(\w[43][31] ),
    .A3(\w[47][31] ),
    .S0(net459),
    .S1(net470),
    .X(_05404_));
 sky130_fd_sc_hd__mux4_2 _15989_ (.A0(\w[49][31] ),
    .A1(\w[53][31] ),
    .A2(\w[51][31] ),
    .A3(\w[55][31] ),
    .S0(net459),
    .S1(net470),
    .X(_05405_));
 sky130_fd_sc_hd__mux4_2 _15990_ (.A0(\w[57][31] ),
    .A1(\w[61][31] ),
    .A2(\w[59][31] ),
    .A3(\w[63][31] ),
    .S0(net459),
    .S1(net470),
    .X(_05406_));
 sky130_fd_sc_hd__mux4_2 _15991_ (.A0(_05403_),
    .A1(_05404_),
    .A2(_05405_),
    .A3(_05406_),
    .S0(net456),
    .S1(net454),
    .X(_05407_));
 sky130_fd_sc_hd__mux2i_4 _15992_ (.A0(_05402_),
    .A1(_05407_),
    .S(net453),
    .Y(_05408_));
 sky130_fd_sc_hd__xnor2_1 _15993_ (.A(_05397_),
    .B(_05408_),
    .Y(_05409_));
 sky130_fd_sc_hd__mux4_2 _15994_ (.A0(\w[0][31] ),
    .A1(\w[4][31] ),
    .A2(\w[2][31] ),
    .A3(\w[6][31] ),
    .S0(net384),
    .S1(net391),
    .X(_05410_));
 sky130_fd_sc_hd__mux4_2 _15995_ (.A0(\w[8][31] ),
    .A1(\w[12][31] ),
    .A2(\w[10][31] ),
    .A3(\w[14][31] ),
    .S0(net384),
    .S1(net391),
    .X(_05411_));
 sky130_fd_sc_hd__mux4_2 _15996_ (.A0(\w[16][31] ),
    .A1(\w[20][31] ),
    .A2(\w[18][31] ),
    .A3(\w[22][31] ),
    .S0(net384),
    .S1(net391),
    .X(_05412_));
 sky130_fd_sc_hd__mux4_2 _15997_ (.A0(\w[24][31] ),
    .A1(\w[28][31] ),
    .A2(\w[26][31] ),
    .A3(\w[30][31] ),
    .S0(net384),
    .S1(net391),
    .X(_05413_));
 sky130_fd_sc_hd__mux4_2 _15998_ (.A0(_05410_),
    .A1(_05411_),
    .A2(_05412_),
    .A3(_05413_),
    .S0(net377),
    .S1(net375),
    .X(_05414_));
 sky130_fd_sc_hd__mux4_2 _15999_ (.A0(\w[32][31] ),
    .A1(\w[36][31] ),
    .A2(\w[34][31] ),
    .A3(\w[38][31] ),
    .S0(net383),
    .S1(net390),
    .X(_05415_));
 sky130_fd_sc_hd__mux4_2 _16000_ (.A0(\w[40][31] ),
    .A1(\w[44][31] ),
    .A2(\w[42][31] ),
    .A3(\w[46][31] ),
    .S0(net383),
    .S1(net390),
    .X(_05416_));
 sky130_fd_sc_hd__mux4_2 _16001_ (.A0(\w[48][31] ),
    .A1(\w[52][31] ),
    .A2(\w[50][31] ),
    .A3(\w[54][31] ),
    .S0(net383),
    .S1(net390),
    .X(_05417_));
 sky130_fd_sc_hd__mux4_2 _16002_ (.A0(\w[56][31] ),
    .A1(\w[60][31] ),
    .A2(\w[58][31] ),
    .A3(\w[62][31] ),
    .S0(net385),
    .S1(net392),
    .X(_05418_));
 sky130_fd_sc_hd__mux4_2 _16003_ (.A0(_05415_),
    .A1(_05416_),
    .A2(_05417_),
    .A3(_05418_),
    .S0(net377),
    .S1(net375),
    .X(_05419_));
 sky130_fd_sc_hd__mux2i_4 _16004_ (.A0(_05414_),
    .A1(_05419_),
    .S(net373),
    .Y(_05420_));
 sky130_fd_sc_hd__xnor2_4 _16005_ (.A(_03656_),
    .B(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__xnor2_1 _16006_ (.A(_05409_),
    .B(_05421_),
    .Y(_05422_));
 sky130_fd_sc_hd__xor2_1 _16007_ (.A(_03194_),
    .B(_03378_),
    .X(_05423_));
 sky130_fd_sc_hd__xnor2_1 _16008_ (.A(_02964_),
    .B(_05423_),
    .Y(_05424_));
 sky130_fd_sc_hd__xnor2_1 _16009_ (.A(_05422_),
    .B(_05424_),
    .Y(_05425_));
 sky130_fd_sc_hd__nor2_1 _16010_ (.A(net351),
    .B(_05425_),
    .Y(_05426_));
 sky130_fd_sc_hd__nand2_1 _16011_ (.A(net339),
    .B(_05425_),
    .Y(_05427_));
 sky130_fd_sc_hd__a21oi_1 _16012_ (.A1(_05393_),
    .A2(_05396_),
    .B1(_05427_),
    .Y(_05428_));
 sky130_fd_sc_hd__nor2_1 _16013_ (.A(\w[63][31] ),
    .B(net339),
    .Y(_05429_));
 sky130_fd_sc_hd__a311o_2 _16014_ (.A1(_05393_),
    .A2(_05396_),
    .A3(_05426_),
    .B1(_05428_),
    .C1(_05429_),
    .X(_05430_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1304 ();
 sky130_fd_sc_hd__nand2_1 _16016_ (.A(net256),
    .B(_05116_),
    .Y(_05432_));
 sky130_fd_sc_hd__o21ai_0 _16017_ (.A1(_05116_),
    .A2(_05430_),
    .B1(_05432_),
    .Y(_00377_));
 sky130_fd_sc_hd__nor2b_4 _16018_ (.A(net1039),
    .B_N(_13531_),
    .Y(_05433_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1303 ();
 sky130_fd_sc_hd__nand2_8 _16020_ (.A(_09735_),
    .B(_05433_),
    .Y(_05435_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1301 ();
 sky130_fd_sc_hd__nand2_1 _16023_ (.A(net774),
    .B(_05435_),
    .Y(_05438_));
 sky130_fd_sc_hd__o21ai_0 _16024_ (.A1(_04790_),
    .A2(_05435_),
    .B1(_05438_),
    .Y(_00385_));
 sky130_fd_sc_hd__nand2_1 _16025_ (.A(net773),
    .B(_05435_),
    .Y(_05439_));
 sky130_fd_sc_hd__o21ai_0 _16026_ (.A1(_04794_),
    .A2(_05435_),
    .B1(_05439_),
    .Y(_00396_));
 sky130_fd_sc_hd__nand2_1 _16027_ (.A(net772),
    .B(_05435_),
    .Y(_05440_));
 sky130_fd_sc_hd__o21ai_0 _16028_ (.A1(_04801_),
    .A2(_05435_),
    .B1(_05440_),
    .Y(_00407_));
 sky130_fd_sc_hd__nand2_1 _16029_ (.A(net771),
    .B(_05435_),
    .Y(_05441_));
 sky130_fd_sc_hd__o21ai_0 _16030_ (.A1(_04808_),
    .A2(_05435_),
    .B1(_05441_),
    .Y(_00410_));
 sky130_fd_sc_hd__nand2_1 _16031_ (.A(net770),
    .B(_05435_),
    .Y(_05442_));
 sky130_fd_sc_hd__o21ai_0 _16032_ (.A1(_04817_),
    .A2(_05435_),
    .B1(_05442_),
    .Y(_00411_));
 sky130_fd_sc_hd__nand2_1 _16033_ (.A(net769),
    .B(_05435_),
    .Y(_05443_));
 sky130_fd_sc_hd__o21ai_0 _16034_ (.A1(_04826_),
    .A2(_05435_),
    .B1(_05443_),
    .Y(_00412_));
 sky130_fd_sc_hd__nand2_1 _16035_ (.A(net767),
    .B(_05435_),
    .Y(_05444_));
 sky130_fd_sc_hd__o21ai_0 _16036_ (.A1(_04834_),
    .A2(_05435_),
    .B1(_05444_),
    .Y(_00413_));
 sky130_fd_sc_hd__nand2_1 _16037_ (.A(net766),
    .B(_05435_),
    .Y(_05445_));
 sky130_fd_sc_hd__o21ai_0 _16038_ (.A1(_04843_),
    .A2(_05435_),
    .B1(_05445_),
    .Y(_00414_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1300 ();
 sky130_fd_sc_hd__nand2_1 _16040_ (.A(net765),
    .B(_05435_),
    .Y(_05447_));
 sky130_fd_sc_hd__o21ai_0 _16041_ (.A1(_04852_),
    .A2(_05435_),
    .B1(_05447_),
    .Y(_00415_));
 sky130_fd_sc_hd__nand2_1 _16042_ (.A(net764),
    .B(_05435_),
    .Y(_05448_));
 sky130_fd_sc_hd__o21ai_0 _16043_ (.A1(_04860_),
    .A2(_05435_),
    .B1(_05448_),
    .Y(_00416_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1299 ();
 sky130_fd_sc_hd__nand2_1 _16045_ (.A(net763),
    .B(_05435_),
    .Y(_05450_));
 sky130_fd_sc_hd__o21ai_0 _16046_ (.A1(_04871_),
    .A2(_05435_),
    .B1(_05450_),
    .Y(_00386_));
 sky130_fd_sc_hd__nand2_1 _16047_ (.A(net762),
    .B(_05435_),
    .Y(_05451_));
 sky130_fd_sc_hd__o21ai_0 _16048_ (.A1(_04883_),
    .A2(_05435_),
    .B1(_05451_),
    .Y(_00387_));
 sky130_fd_sc_hd__nand2_1 _16049_ (.A(net761),
    .B(_05435_),
    .Y(_05452_));
 sky130_fd_sc_hd__o21ai_0 _16050_ (.A1(_04892_),
    .A2(_05435_),
    .B1(_05452_),
    .Y(_00388_));
 sky130_fd_sc_hd__nand2_1 _16051_ (.A(net760),
    .B(_05435_),
    .Y(_05453_));
 sky130_fd_sc_hd__o21ai_0 _16052_ (.A1(_04899_),
    .A2(_05435_),
    .B1(_05453_),
    .Y(_00389_));
 sky130_fd_sc_hd__nand2_1 _16053_ (.A(net759),
    .B(_05435_),
    .Y(_05454_));
 sky130_fd_sc_hd__o21ai_0 _16054_ (.A1(_04906_),
    .A2(_05435_),
    .B1(_05454_),
    .Y(_00390_));
 sky130_fd_sc_hd__nand2_1 _16055_ (.A(net758),
    .B(_05435_),
    .Y(_05455_));
 sky130_fd_sc_hd__o21ai_0 _16056_ (.A1(_04913_),
    .A2(_05435_),
    .B1(_05455_),
    .Y(_00391_));
 sky130_fd_sc_hd__nand2_1 _16057_ (.A(net756),
    .B(_05435_),
    .Y(_05456_));
 sky130_fd_sc_hd__o21ai_0 _16058_ (.A1(_04923_),
    .A2(_05435_),
    .B1(_05456_),
    .Y(_00392_));
 sky130_fd_sc_hd__nand2_1 _16059_ (.A(net755),
    .B(_05435_),
    .Y(_05457_));
 sky130_fd_sc_hd__o21ai_0 _16060_ (.A1(_04932_),
    .A2(_05435_),
    .B1(_05457_),
    .Y(_00393_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1298 ();
 sky130_fd_sc_hd__nand2_1 _16062_ (.A(net754),
    .B(_05435_),
    .Y(_05459_));
 sky130_fd_sc_hd__o21ai_0 _16063_ (.A1(_04939_),
    .A2(_05435_),
    .B1(_05459_),
    .Y(_00394_));
 sky130_fd_sc_hd__nand2_1 _16064_ (.A(net753),
    .B(_05435_),
    .Y(_05460_));
 sky130_fd_sc_hd__o21ai_0 _16065_ (.A1(_04951_),
    .A2(_05435_),
    .B1(_05460_),
    .Y(_00395_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1297 ();
 sky130_fd_sc_hd__nand2_1 _16067_ (.A(net752),
    .B(_05435_),
    .Y(_05462_));
 sky130_fd_sc_hd__o21ai_0 _16068_ (.A1(_04960_),
    .A2(_05435_),
    .B1(_05462_),
    .Y(_00397_));
 sky130_fd_sc_hd__nand2_1 _16069_ (.A(net751),
    .B(_05435_),
    .Y(_05463_));
 sky130_fd_sc_hd__o21ai_0 _16070_ (.A1(_04974_),
    .A2(_05435_),
    .B1(_05463_),
    .Y(_00398_));
 sky130_fd_sc_hd__nand2_1 _16071_ (.A(net750),
    .B(_05435_),
    .Y(_05464_));
 sky130_fd_sc_hd__o21ai_0 _16072_ (.A1(_04984_),
    .A2(_05435_),
    .B1(_05464_),
    .Y(_00399_));
 sky130_fd_sc_hd__nand2_1 _16073_ (.A(net749),
    .B(_05435_),
    .Y(_05465_));
 sky130_fd_sc_hd__o21ai_0 _16074_ (.A1(_04990_),
    .A2(_05435_),
    .B1(_05465_),
    .Y(_00400_));
 sky130_fd_sc_hd__nand2_1 _16075_ (.A(net748),
    .B(_05435_),
    .Y(_05466_));
 sky130_fd_sc_hd__o21ai_0 _16076_ (.A1(net1129),
    .A2(_05435_),
    .B1(_05466_),
    .Y(_00401_));
 sky130_fd_sc_hd__nand2_1 _16077_ (.A(net747),
    .B(_05435_),
    .Y(_05467_));
 sky130_fd_sc_hd__o21ai_0 _16078_ (.A1(_05011_),
    .A2(_05435_),
    .B1(_05467_),
    .Y(_00402_));
 sky130_fd_sc_hd__nand2_1 _16079_ (.A(net745),
    .B(_05435_),
    .Y(_05468_));
 sky130_fd_sc_hd__o21ai_0 _16080_ (.A1(_05020_),
    .A2(_05435_),
    .B1(_05468_),
    .Y(_00403_));
 sky130_fd_sc_hd__nand2_1 _16081_ (.A(net744),
    .B(_05435_),
    .Y(_05469_));
 sky130_fd_sc_hd__o21ai_0 _16082_ (.A1(_05029_),
    .A2(_05435_),
    .B1(_05469_),
    .Y(_00404_));
 sky130_fd_sc_hd__nand2_1 _16083_ (.A(net743),
    .B(_05435_),
    .Y(_05470_));
 sky130_fd_sc_hd__o21ai_0 _16084_ (.A1(_05035_),
    .A2(_05435_),
    .B1(_05470_),
    .Y(_00405_));
 sky130_fd_sc_hd__nand2_1 _16085_ (.A(net742),
    .B(_05435_),
    .Y(_05471_));
 sky130_fd_sc_hd__o21ai_0 _16086_ (.A1(_05044_),
    .A2(_05435_),
    .B1(_05471_),
    .Y(_00406_));
 sky130_fd_sc_hd__nand2_1 _16087_ (.A(net741),
    .B(_05435_),
    .Y(_05472_));
 sky130_fd_sc_hd__o21ai_0 _16088_ (.A1(_05060_),
    .A2(_05435_),
    .B1(_05472_),
    .Y(_00408_));
 sky130_fd_sc_hd__mux2i_1 _16089_ (.A0(_05113_),
    .A1(net740),
    .S(_05435_),
    .Y(_05473_));
 sky130_fd_sc_hd__o21ai_0 _16090_ (.A1(_05112_),
    .A2(_05435_),
    .B1(_05473_),
    .Y(_00409_));
 sky130_fd_sc_hd__nor2b_4 _16091_ (.A(net1039),
    .B_N(_13539_),
    .Y(_05474_));
 sky130_fd_sc_hd__nand2_8 _16092_ (.A(_09797_),
    .B(_05474_),
    .Y(_05475_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1295 ();
 sky130_fd_sc_hd__nand2_1 _16095_ (.A(net31),
    .B(_05475_),
    .Y(_05478_));
 sky130_fd_sc_hd__o21ai_0 _16096_ (.A1(_05118_),
    .A2(_05475_),
    .B1(_05478_),
    .Y(_00417_));
 sky130_fd_sc_hd__nand2_1 _16097_ (.A(net30),
    .B(_05475_),
    .Y(_05479_));
 sky130_fd_sc_hd__o21ai_0 _16098_ (.A1(_05122_),
    .A2(_05475_),
    .B1(_05479_),
    .Y(_00428_));
 sky130_fd_sc_hd__nand2_1 _16099_ (.A(net29),
    .B(_05475_),
    .Y(_05480_));
 sky130_fd_sc_hd__o21ai_0 _16100_ (.A1(_05126_),
    .A2(_05475_),
    .B1(_05480_),
    .Y(_00439_));
 sky130_fd_sc_hd__nand2_1 _16101_ (.A(net28),
    .B(_05475_),
    .Y(_05481_));
 sky130_fd_sc_hd__o21ai_0 _16102_ (.A1(_05132_),
    .A2(_05475_),
    .B1(_05481_),
    .Y(_00442_));
 sky130_fd_sc_hd__nand2_1 _16103_ (.A(net27),
    .B(_05475_),
    .Y(_05482_));
 sky130_fd_sc_hd__o21ai_0 _16104_ (.A1(_05140_),
    .A2(_05475_),
    .B1(_05482_),
    .Y(_00443_));
 sky130_fd_sc_hd__nand2_1 _16105_ (.A(net26),
    .B(_05475_),
    .Y(_05483_));
 sky130_fd_sc_hd__o21ai_0 _16106_ (.A1(_05149_),
    .A2(_05475_),
    .B1(_05483_),
    .Y(_00444_));
 sky130_fd_sc_hd__nand2_1 _16107_ (.A(net25),
    .B(_05475_),
    .Y(_05484_));
 sky130_fd_sc_hd__o21ai_0 _16108_ (.A1(_05157_),
    .A2(_05475_),
    .B1(_05484_),
    .Y(_00445_));
 sky130_fd_sc_hd__nand2_1 _16109_ (.A(net24),
    .B(_05475_),
    .Y(_05485_));
 sky130_fd_sc_hd__o21ai_0 _16110_ (.A1(_05166_),
    .A2(_05475_),
    .B1(_05485_),
    .Y(_00446_));
 sky130_fd_sc_hd__nand2_1 _16111_ (.A(net22),
    .B(_05475_),
    .Y(_05486_));
 sky130_fd_sc_hd__o21ai_0 _16112_ (.A1(_05173_),
    .A2(_05475_),
    .B1(_05486_),
    .Y(_00447_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1294 ();
 sky130_fd_sc_hd__nand2_1 _16114_ (.A(net21),
    .B(_05475_),
    .Y(_05488_));
 sky130_fd_sc_hd__o21ai_0 _16115_ (.A1(_05183_),
    .A2(_05475_),
    .B1(_05488_),
    .Y(_00448_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1293 ();
 sky130_fd_sc_hd__nand2_1 _16117_ (.A(net20),
    .B(_05475_),
    .Y(_05490_));
 sky130_fd_sc_hd__o21ai_0 _16118_ (.A1(_05192_),
    .A2(_05475_),
    .B1(_05490_),
    .Y(_00418_));
 sky130_fd_sc_hd__nand2_1 _16119_ (.A(net19),
    .B(_05475_),
    .Y(_05491_));
 sky130_fd_sc_hd__o21ai_0 _16120_ (.A1(_05204_),
    .A2(_05475_),
    .B1(_05491_),
    .Y(_00419_));
 sky130_fd_sc_hd__nand2_1 _16121_ (.A(net18),
    .B(_05475_),
    .Y(_05492_));
 sky130_fd_sc_hd__o21ai_0 _16122_ (.A1(_05214_),
    .A2(_05475_),
    .B1(_05492_),
    .Y(_00420_));
 sky130_fd_sc_hd__nand2_1 _16123_ (.A(net17),
    .B(_05475_),
    .Y(_05493_));
 sky130_fd_sc_hd__o21ai_0 _16124_ (.A1(_05221_),
    .A2(_05475_),
    .B1(_05493_),
    .Y(_00421_));
 sky130_fd_sc_hd__nand2_1 _16125_ (.A(net16),
    .B(_05475_),
    .Y(_05494_));
 sky130_fd_sc_hd__o21ai_0 _16126_ (.A1(_05228_),
    .A2(_05475_),
    .B1(_05494_),
    .Y(_00422_));
 sky130_fd_sc_hd__nand2_1 _16127_ (.A(net15),
    .B(_05475_),
    .Y(_05495_));
 sky130_fd_sc_hd__o21ai_0 _16128_ (.A1(_05238_),
    .A2(_05475_),
    .B1(_05495_),
    .Y(_00423_));
 sky130_fd_sc_hd__nand2_1 _16129_ (.A(net14),
    .B(_05475_),
    .Y(_05496_));
 sky130_fd_sc_hd__o21ai_0 _16130_ (.A1(_05247_),
    .A2(_05475_),
    .B1(_05496_),
    .Y(_00424_));
 sky130_fd_sc_hd__nand2_1 _16131_ (.A(net13),
    .B(_05475_),
    .Y(_05497_));
 sky130_fd_sc_hd__o21ai_0 _16132_ (.A1(_05258_),
    .A2(_05475_),
    .B1(_05497_),
    .Y(_00425_));
 sky130_fd_sc_hd__nand2_1 _16133_ (.A(net11),
    .B(_05475_),
    .Y(_05498_));
 sky130_fd_sc_hd__o21ai_0 _16134_ (.A1(_05267_),
    .A2(_05475_),
    .B1(_05498_),
    .Y(_00426_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1292 ();
 sky130_fd_sc_hd__nand2_1 _16136_ (.A(net10),
    .B(_05475_),
    .Y(_05500_));
 sky130_fd_sc_hd__o21ai_0 _16137_ (.A1(_05280_),
    .A2(_05475_),
    .B1(_05500_),
    .Y(_00427_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1291 ();
 sky130_fd_sc_hd__nand2_1 _16139_ (.A(net9),
    .B(_05475_),
    .Y(_05502_));
 sky130_fd_sc_hd__o21ai_0 _16140_ (.A1(_05291_),
    .A2(_05475_),
    .B1(_05502_),
    .Y(_00429_));
 sky130_fd_sc_hd__nand2_1 _16141_ (.A(net8),
    .B(_05475_),
    .Y(_05503_));
 sky130_fd_sc_hd__o21ai_0 _16142_ (.A1(_05301_),
    .A2(_05475_),
    .B1(_05503_),
    .Y(_00430_));
 sky130_fd_sc_hd__nand2_1 _16143_ (.A(net7),
    .B(_05475_),
    .Y(_05504_));
 sky130_fd_sc_hd__o21ai_0 _16144_ (.A1(_05309_),
    .A2(_05475_),
    .B1(_05504_),
    .Y(_00431_));
 sky130_fd_sc_hd__nand2_1 _16145_ (.A(net6),
    .B(_05475_),
    .Y(_05505_));
 sky130_fd_sc_hd__o21ai_0 _16146_ (.A1(_05320_),
    .A2(_05475_),
    .B1(_05505_),
    .Y(_00432_));
 sky130_fd_sc_hd__nand2_1 _16147_ (.A(net5),
    .B(_05475_),
    .Y(_05506_));
 sky130_fd_sc_hd__o21ai_0 _16148_ (.A1(net1145),
    .A2(_05475_),
    .B1(_05506_),
    .Y(_00433_));
 sky130_fd_sc_hd__nand2_1 _16149_ (.A(net4),
    .B(_05475_),
    .Y(_05507_));
 sky130_fd_sc_hd__o21ai_0 _16150_ (.A1(_05339_),
    .A2(_05475_),
    .B1(_05507_),
    .Y(_00434_));
 sky130_fd_sc_hd__nand2_1 _16151_ (.A(net3),
    .B(_05475_),
    .Y(_05508_));
 sky130_fd_sc_hd__o21ai_0 _16152_ (.A1(_05347_),
    .A2(_05475_),
    .B1(_05508_),
    .Y(_00435_));
 sky130_fd_sc_hd__nand2_1 _16153_ (.A(net2),
    .B(_05475_),
    .Y(_05509_));
 sky130_fd_sc_hd__o21ai_0 _16154_ (.A1(_05358_),
    .A2(_05475_),
    .B1(_05509_),
    .Y(_00436_));
 sky130_fd_sc_hd__nand2_1 _16155_ (.A(net778),
    .B(_05475_),
    .Y(_05510_));
 sky130_fd_sc_hd__o21ai_0 _16156_ (.A1(_05372_),
    .A2(_05475_),
    .B1(_05510_),
    .Y(_00437_));
 sky130_fd_sc_hd__nand2_1 _16157_ (.A(net777),
    .B(_05475_),
    .Y(_05511_));
 sky130_fd_sc_hd__o21ai_0 _16158_ (.A1(_05380_),
    .A2(_05475_),
    .B1(_05511_),
    .Y(_00438_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1289 ();
 sky130_fd_sc_hd__a21oi_1 _16161_ (.A1(_09797_),
    .A2(_05474_),
    .B1(net776),
    .Y(_05514_));
 sky130_fd_sc_hd__a31oi_1 _16162_ (.A1(_09797_),
    .A2(net1143),
    .A3(_05474_),
    .B1(_05514_),
    .Y(_00440_));
 sky130_fd_sc_hd__nand2_1 _16163_ (.A(net775),
    .B(_05475_),
    .Y(_05515_));
 sky130_fd_sc_hd__o21ai_0 _16164_ (.A1(_05430_),
    .A2(_05475_),
    .B1(_05515_),
    .Y(_00441_));
 sky130_fd_sc_hd__nor2b_4 _16165_ (.A(net1038),
    .B_N(_13529_),
    .Y(_05516_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1288 ();
 sky130_fd_sc_hd__nand2_8 _16167_ (.A(_09735_),
    .B(_05516_),
    .Y(_05518_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1286 ();
 sky130_fd_sc_hd__nand2_1 _16170_ (.A(net66),
    .B(_05518_),
    .Y(_05521_));
 sky130_fd_sc_hd__o21ai_0 _16171_ (.A1(_04790_),
    .A2(_05518_),
    .B1(_05521_),
    .Y(_00449_));
 sky130_fd_sc_hd__nand2_1 _16172_ (.A(net65),
    .B(_05518_),
    .Y(_05522_));
 sky130_fd_sc_hd__o21ai_0 _16173_ (.A1(_04794_),
    .A2(_05518_),
    .B1(_05522_),
    .Y(_00460_));
 sky130_fd_sc_hd__nand2_1 _16174_ (.A(net64),
    .B(_05518_),
    .Y(_05523_));
 sky130_fd_sc_hd__o21ai_0 _16175_ (.A1(_04801_),
    .A2(_05518_),
    .B1(_05523_),
    .Y(_00471_));
 sky130_fd_sc_hd__nand2_1 _16176_ (.A(net63),
    .B(_05518_),
    .Y(_05524_));
 sky130_fd_sc_hd__o21ai_0 _16177_ (.A1(_04808_),
    .A2(_05518_),
    .B1(_05524_),
    .Y(_00474_));
 sky130_fd_sc_hd__nand2_1 _16178_ (.A(net62),
    .B(_05518_),
    .Y(_05525_));
 sky130_fd_sc_hd__o21ai_0 _16179_ (.A1(_04817_),
    .A2(_05518_),
    .B1(_05525_),
    .Y(_00475_));
 sky130_fd_sc_hd__nand2_1 _16180_ (.A(net61),
    .B(_05518_),
    .Y(_05526_));
 sky130_fd_sc_hd__o21ai_0 _16181_ (.A1(_04826_),
    .A2(_05518_),
    .B1(_05526_),
    .Y(_00476_));
 sky130_fd_sc_hd__nand2_1 _16182_ (.A(net60),
    .B(_05518_),
    .Y(_05527_));
 sky130_fd_sc_hd__o21ai_0 _16183_ (.A1(_04834_),
    .A2(_05518_),
    .B1(_05527_),
    .Y(_00477_));
 sky130_fd_sc_hd__nand2_1 _16184_ (.A(net59),
    .B(_05518_),
    .Y(_05528_));
 sky130_fd_sc_hd__o21ai_0 _16185_ (.A1(_04843_),
    .A2(_05518_),
    .B1(_05528_),
    .Y(_00478_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1285 ();
 sky130_fd_sc_hd__nand2_1 _16187_ (.A(net58),
    .B(_05518_),
    .Y(_05530_));
 sky130_fd_sc_hd__o21ai_0 _16188_ (.A1(_04852_),
    .A2(_05518_),
    .B1(_05530_),
    .Y(_00479_));
 sky130_fd_sc_hd__nand2_1 _16189_ (.A(net57),
    .B(_05518_),
    .Y(_05531_));
 sky130_fd_sc_hd__o21ai_0 _16190_ (.A1(_04860_),
    .A2(_05518_),
    .B1(_05531_),
    .Y(_00480_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1284 ();
 sky130_fd_sc_hd__nand2_1 _16192_ (.A(net55),
    .B(_05518_),
    .Y(_05533_));
 sky130_fd_sc_hd__o21ai_0 _16193_ (.A1(_04871_),
    .A2(_05518_),
    .B1(_05533_),
    .Y(_00450_));
 sky130_fd_sc_hd__nand2_1 _16194_ (.A(net54),
    .B(_05518_),
    .Y(_05534_));
 sky130_fd_sc_hd__o21ai_0 _16195_ (.A1(_04883_),
    .A2(_05518_),
    .B1(_05534_),
    .Y(_00451_));
 sky130_fd_sc_hd__nand2_1 _16196_ (.A(net53),
    .B(_05518_),
    .Y(_05535_));
 sky130_fd_sc_hd__o21ai_0 _16197_ (.A1(_04892_),
    .A2(_05518_),
    .B1(_05535_),
    .Y(_00452_));
 sky130_fd_sc_hd__nand2_1 _16198_ (.A(net52),
    .B(_05518_),
    .Y(_05536_));
 sky130_fd_sc_hd__o21ai_0 _16199_ (.A1(_04899_),
    .A2(_05518_),
    .B1(_05536_),
    .Y(_00453_));
 sky130_fd_sc_hd__nand2_1 _16200_ (.A(net51),
    .B(_05518_),
    .Y(_05537_));
 sky130_fd_sc_hd__o21ai_0 _16201_ (.A1(_04906_),
    .A2(_05518_),
    .B1(_05537_),
    .Y(_00454_));
 sky130_fd_sc_hd__nand2_1 _16202_ (.A(net50),
    .B(_05518_),
    .Y(_05538_));
 sky130_fd_sc_hd__o21ai_0 _16203_ (.A1(_04913_),
    .A2(_05518_),
    .B1(_05538_),
    .Y(_00455_));
 sky130_fd_sc_hd__nand2_1 _16204_ (.A(net49),
    .B(_05518_),
    .Y(_05539_));
 sky130_fd_sc_hd__o21ai_0 _16205_ (.A1(_04923_),
    .A2(_05518_),
    .B1(_05539_),
    .Y(_00456_));
 sky130_fd_sc_hd__nand2_1 _16206_ (.A(net48),
    .B(_05518_),
    .Y(_05540_));
 sky130_fd_sc_hd__o21ai_0 _16207_ (.A1(_04932_),
    .A2(_05518_),
    .B1(_05540_),
    .Y(_00457_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1283 ();
 sky130_fd_sc_hd__nand2_1 _16209_ (.A(net47),
    .B(_05518_),
    .Y(_05542_));
 sky130_fd_sc_hd__o21ai_0 _16210_ (.A1(_04939_),
    .A2(_05518_),
    .B1(_05542_),
    .Y(_00458_));
 sky130_fd_sc_hd__nand2_1 _16211_ (.A(net46),
    .B(_05518_),
    .Y(_05543_));
 sky130_fd_sc_hd__o21ai_0 _16212_ (.A1(_04951_),
    .A2(_05518_),
    .B1(_05543_),
    .Y(_00459_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1282 ();
 sky130_fd_sc_hd__nand2_1 _16214_ (.A(net44),
    .B(_05518_),
    .Y(_05545_));
 sky130_fd_sc_hd__o21ai_0 _16215_ (.A1(_04960_),
    .A2(_05518_),
    .B1(_05545_),
    .Y(_00461_));
 sky130_fd_sc_hd__nand2_1 _16216_ (.A(net43),
    .B(_05518_),
    .Y(_05546_));
 sky130_fd_sc_hd__o21ai_0 _16217_ (.A1(_04974_),
    .A2(_05518_),
    .B1(_05546_),
    .Y(_00462_));
 sky130_fd_sc_hd__nand2_1 _16218_ (.A(net42),
    .B(_05518_),
    .Y(_05547_));
 sky130_fd_sc_hd__o21ai_0 _16219_ (.A1(_04984_),
    .A2(_05518_),
    .B1(_05547_),
    .Y(_00463_));
 sky130_fd_sc_hd__nand2_1 _16220_ (.A(net41),
    .B(_05518_),
    .Y(_05548_));
 sky130_fd_sc_hd__o21ai_0 _16221_ (.A1(_04990_),
    .A2(_05518_),
    .B1(_05548_),
    .Y(_00464_));
 sky130_fd_sc_hd__nand2_1 _16222_ (.A(net40),
    .B(_05518_),
    .Y(_05549_));
 sky130_fd_sc_hd__o21ai_0 _16223_ (.A1(net1129),
    .A2(_05518_),
    .B1(_05549_),
    .Y(_00465_));
 sky130_fd_sc_hd__nand2_1 _16224_ (.A(net39),
    .B(_05518_),
    .Y(_05550_));
 sky130_fd_sc_hd__o21ai_0 _16225_ (.A1(_05011_),
    .A2(_05518_),
    .B1(_05550_),
    .Y(_00466_));
 sky130_fd_sc_hd__nand2_1 _16226_ (.A(net38),
    .B(_05518_),
    .Y(_05551_));
 sky130_fd_sc_hd__o21ai_0 _16227_ (.A1(_05020_),
    .A2(_05518_),
    .B1(_05551_),
    .Y(_00467_));
 sky130_fd_sc_hd__nand2_1 _16228_ (.A(net37),
    .B(_05518_),
    .Y(_05552_));
 sky130_fd_sc_hd__o21ai_0 _16229_ (.A1(_05029_),
    .A2(_05518_),
    .B1(_05552_),
    .Y(_00468_));
 sky130_fd_sc_hd__nand2_1 _16230_ (.A(net36),
    .B(_05518_),
    .Y(_05553_));
 sky130_fd_sc_hd__o21ai_0 _16231_ (.A1(_05035_),
    .A2(_05518_),
    .B1(_05553_),
    .Y(_00469_));
 sky130_fd_sc_hd__nand2_1 _16232_ (.A(net35),
    .B(_05518_),
    .Y(_05554_));
 sky130_fd_sc_hd__o21ai_0 _16233_ (.A1(_05044_),
    .A2(_05518_),
    .B1(_05554_),
    .Y(_00470_));
 sky130_fd_sc_hd__nand2_1 _16234_ (.A(net33),
    .B(_05518_),
    .Y(_05555_));
 sky130_fd_sc_hd__o21ai_0 _16235_ (.A1(_05060_),
    .A2(_05518_),
    .B1(_05555_),
    .Y(_00472_));
 sky130_fd_sc_hd__mux2i_1 _16236_ (.A0(_05113_),
    .A1(net32),
    .S(_05518_),
    .Y(_05556_));
 sky130_fd_sc_hd__o21ai_0 _16237_ (.A1(_05112_),
    .A2(_05518_),
    .B1(_05556_),
    .Y(_00473_));
 sky130_fd_sc_hd__nor2b_4 _16238_ (.A(net1039),
    .B_N(_13537_),
    .Y(_05557_));
 sky130_fd_sc_hd__nand2_8 _16239_ (.A(_09797_),
    .B(_05557_),
    .Y(_05558_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1280 ();
 sky130_fd_sc_hd__nand2_1 _16242_ (.A(net102),
    .B(_05558_),
    .Y(_05561_));
 sky130_fd_sc_hd__o21ai_0 _16243_ (.A1(_05118_),
    .A2(_05558_),
    .B1(_05561_),
    .Y(_00481_));
 sky130_fd_sc_hd__nand2_1 _16244_ (.A(net101),
    .B(_05558_),
    .Y(_05562_));
 sky130_fd_sc_hd__o21ai_0 _16245_ (.A1(_05122_),
    .A2(_05558_),
    .B1(_05562_),
    .Y(_00492_));
 sky130_fd_sc_hd__nand2_1 _16246_ (.A(net99),
    .B(_05558_),
    .Y(_05563_));
 sky130_fd_sc_hd__o21ai_0 _16247_ (.A1(_05126_),
    .A2(_05558_),
    .B1(_05563_),
    .Y(_00503_));
 sky130_fd_sc_hd__nand2_1 _16248_ (.A(net98),
    .B(_05558_),
    .Y(_05564_));
 sky130_fd_sc_hd__o21ai_0 _16249_ (.A1(_05132_),
    .A2(_05558_),
    .B1(_05564_),
    .Y(_00506_));
 sky130_fd_sc_hd__nand2_1 _16250_ (.A(net97),
    .B(_05558_),
    .Y(_05565_));
 sky130_fd_sc_hd__o21ai_0 _16251_ (.A1(_05140_),
    .A2(_05558_),
    .B1(_05565_),
    .Y(_00507_));
 sky130_fd_sc_hd__nand2_1 _16252_ (.A(net96),
    .B(_05558_),
    .Y(_05566_));
 sky130_fd_sc_hd__o21ai_0 _16253_ (.A1(_05149_),
    .A2(_05558_),
    .B1(_05566_),
    .Y(_00508_));
 sky130_fd_sc_hd__nand2_1 _16254_ (.A(net95),
    .B(_05558_),
    .Y(_05567_));
 sky130_fd_sc_hd__o21ai_0 _16255_ (.A1(_05157_),
    .A2(_05558_),
    .B1(_05567_),
    .Y(_00509_));
 sky130_fd_sc_hd__nand2_2 _16256_ (.A(net94),
    .B(_05558_),
    .Y(_05568_));
 sky130_fd_sc_hd__o21ai_0 _16257_ (.A1(_05166_),
    .A2(_05558_),
    .B1(_05568_),
    .Y(_00510_));
 sky130_fd_sc_hd__nand2_1 _16258_ (.A(net93),
    .B(_05558_),
    .Y(_05569_));
 sky130_fd_sc_hd__o21ai_0 _16259_ (.A1(_05173_),
    .A2(_05558_),
    .B1(_05569_),
    .Y(_00511_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1279 ();
 sky130_fd_sc_hd__nand2_1 _16261_ (.A(net92),
    .B(_05558_),
    .Y(_05571_));
 sky130_fd_sc_hd__o21ai_0 _16262_ (.A1(_05183_),
    .A2(_05558_),
    .B1(_05571_),
    .Y(_00512_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1278 ();
 sky130_fd_sc_hd__nand2_1 _16264_ (.A(net91),
    .B(_05558_),
    .Y(_05573_));
 sky130_fd_sc_hd__o21ai_0 _16265_ (.A1(_05192_),
    .A2(_05558_),
    .B1(_05573_),
    .Y(_00482_));
 sky130_fd_sc_hd__nand2_1 _16266_ (.A(net90),
    .B(_05558_),
    .Y(_05574_));
 sky130_fd_sc_hd__o21ai_0 _16267_ (.A1(_05204_),
    .A2(_05558_),
    .B1(_05574_),
    .Y(_00483_));
 sky130_fd_sc_hd__nand2_1 _16268_ (.A(net88),
    .B(_05558_),
    .Y(_05575_));
 sky130_fd_sc_hd__o21ai_0 _16269_ (.A1(_05214_),
    .A2(_05558_),
    .B1(_05575_),
    .Y(_00484_));
 sky130_fd_sc_hd__nand2_1 _16270_ (.A(net87),
    .B(_05558_),
    .Y(_05576_));
 sky130_fd_sc_hd__o21ai_0 _16271_ (.A1(_05221_),
    .A2(_05558_),
    .B1(_05576_),
    .Y(_00485_));
 sky130_fd_sc_hd__nand2_1 _16272_ (.A(net86),
    .B(_05558_),
    .Y(_05577_));
 sky130_fd_sc_hd__o21ai_0 _16273_ (.A1(_05228_),
    .A2(_05558_),
    .B1(_05577_),
    .Y(_00486_));
 sky130_fd_sc_hd__nand2_1 _16274_ (.A(net85),
    .B(_05558_),
    .Y(_05578_));
 sky130_fd_sc_hd__o21ai_0 _16275_ (.A1(_05238_),
    .A2(_05558_),
    .B1(_05578_),
    .Y(_00487_));
 sky130_fd_sc_hd__nand2_1 _16276_ (.A(net84),
    .B(_05558_),
    .Y(_05579_));
 sky130_fd_sc_hd__o21ai_0 _16277_ (.A1(_05247_),
    .A2(_05558_),
    .B1(_05579_),
    .Y(_00488_));
 sky130_fd_sc_hd__nand2_1 _16278_ (.A(net83),
    .B(_05558_),
    .Y(_05580_));
 sky130_fd_sc_hd__o21ai_0 _16279_ (.A1(_05258_),
    .A2(_05558_),
    .B1(_05580_),
    .Y(_00489_));
 sky130_fd_sc_hd__nand2_1 _16280_ (.A(net82),
    .B(_05558_),
    .Y(_05581_));
 sky130_fd_sc_hd__o21ai_0 _16281_ (.A1(_05267_),
    .A2(_05558_),
    .B1(_05581_),
    .Y(_00490_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1277 ();
 sky130_fd_sc_hd__nand2_1 _16283_ (.A(net81),
    .B(_05558_),
    .Y(_05583_));
 sky130_fd_sc_hd__o21ai_0 _16284_ (.A1(_05280_),
    .A2(_05558_),
    .B1(_05583_),
    .Y(_00491_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1276 ();
 sky130_fd_sc_hd__nand2_1 _16286_ (.A(net80),
    .B(_05558_),
    .Y(_05585_));
 sky130_fd_sc_hd__o21ai_0 _16287_ (.A1(_05291_),
    .A2(_05558_),
    .B1(_05585_),
    .Y(_00493_));
 sky130_fd_sc_hd__nand2_1 _16288_ (.A(net79),
    .B(_05558_),
    .Y(_05586_));
 sky130_fd_sc_hd__o21ai_0 _16289_ (.A1(_05301_),
    .A2(_05558_),
    .B1(_05586_),
    .Y(_00494_));
 sky130_fd_sc_hd__nand2_1 _16290_ (.A(net77),
    .B(_05558_),
    .Y(_05587_));
 sky130_fd_sc_hd__o21ai_0 _16291_ (.A1(_05309_),
    .A2(_05558_),
    .B1(_05587_),
    .Y(_00495_));
 sky130_fd_sc_hd__nand2_1 _16292_ (.A(net76),
    .B(_05558_),
    .Y(_05588_));
 sky130_fd_sc_hd__o21ai_0 _16293_ (.A1(_05320_),
    .A2(_05558_),
    .B1(_05588_),
    .Y(_00496_));
 sky130_fd_sc_hd__nand2_1 _16294_ (.A(net75),
    .B(_05558_),
    .Y(_05589_));
 sky130_fd_sc_hd__o21ai_0 _16295_ (.A1(net1145),
    .A2(_05558_),
    .B1(_05589_),
    .Y(_00497_));
 sky130_fd_sc_hd__nand2_1 _16296_ (.A(net74),
    .B(_05558_),
    .Y(_05590_));
 sky130_fd_sc_hd__o21ai_0 _16297_ (.A1(_05339_),
    .A2(_05558_),
    .B1(_05590_),
    .Y(_00498_));
 sky130_fd_sc_hd__nand2_1 _16298_ (.A(net73),
    .B(_05558_),
    .Y(_05591_));
 sky130_fd_sc_hd__o21ai_0 _16299_ (.A1(_05347_),
    .A2(_05558_),
    .B1(_05591_),
    .Y(_00499_));
 sky130_fd_sc_hd__nand2_1 _16300_ (.A(net72),
    .B(_05558_),
    .Y(_05592_));
 sky130_fd_sc_hd__o21ai_0 _16301_ (.A1(_05358_),
    .A2(_05558_),
    .B1(_05592_),
    .Y(_00500_));
 sky130_fd_sc_hd__nand2_1 _16302_ (.A(net71),
    .B(_05558_),
    .Y(_05593_));
 sky130_fd_sc_hd__o21ai_0 _16303_ (.A1(_05372_),
    .A2(_05558_),
    .B1(_05593_),
    .Y(_00501_));
 sky130_fd_sc_hd__nand2_1 _16304_ (.A(net70),
    .B(_05558_),
    .Y(_05594_));
 sky130_fd_sc_hd__o21ai_0 _16305_ (.A1(_05380_),
    .A2(_05558_),
    .B1(_05594_),
    .Y(_00502_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1275 ();
 sky130_fd_sc_hd__a21oi_1 _16307_ (.A1(_09797_),
    .A2(_05557_),
    .B1(net69),
    .Y(_05596_));
 sky130_fd_sc_hd__a31oi_1 _16308_ (.A1(_09797_),
    .A2(net1143),
    .A3(_05557_),
    .B1(_05596_),
    .Y(_00504_));
 sky130_fd_sc_hd__nand2_1 _16309_ (.A(net68),
    .B(_05558_),
    .Y(_05597_));
 sky130_fd_sc_hd__o21ai_0 _16310_ (.A1(_05430_),
    .A2(_05558_),
    .B1(_05597_),
    .Y(_00505_));
 sky130_fd_sc_hd__nor2b_4 _16311_ (.A(net1039),
    .B_N(_13533_),
    .Y(_05598_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1274 ();
 sky130_fd_sc_hd__nand2_8 _16313_ (.A(_09735_),
    .B(_05598_),
    .Y(_05600_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1272 ();
 sky130_fd_sc_hd__nand2_1 _16316_ (.A(net138),
    .B(_05600_),
    .Y(_05603_));
 sky130_fd_sc_hd__o21ai_0 _16317_ (.A1(_04790_),
    .A2(_05600_),
    .B1(_05603_),
    .Y(_00513_));
 sky130_fd_sc_hd__nand2_1 _16318_ (.A(net137),
    .B(_05600_),
    .Y(_05604_));
 sky130_fd_sc_hd__o21ai_0 _16319_ (.A1(_04794_),
    .A2(_05600_),
    .B1(_05604_),
    .Y(_00524_));
 sky130_fd_sc_hd__nand2_1 _16320_ (.A(net136),
    .B(_05600_),
    .Y(_05605_));
 sky130_fd_sc_hd__o21ai_0 _16321_ (.A1(_04801_),
    .A2(_05600_),
    .B1(_05605_),
    .Y(_00535_));
 sky130_fd_sc_hd__nand2_1 _16322_ (.A(net135),
    .B(_05600_),
    .Y(_05606_));
 sky130_fd_sc_hd__o21ai_0 _16323_ (.A1(_04808_),
    .A2(_05600_),
    .B1(_05606_),
    .Y(_00538_));
 sky130_fd_sc_hd__nand2_1 _16324_ (.A(net133),
    .B(_05600_),
    .Y(_05607_));
 sky130_fd_sc_hd__o21ai_0 _16325_ (.A1(_04817_),
    .A2(_05600_),
    .B1(_05607_),
    .Y(_00539_));
 sky130_fd_sc_hd__nand2_1 _16326_ (.A(net132),
    .B(_05600_),
    .Y(_05608_));
 sky130_fd_sc_hd__o21ai_0 _16327_ (.A1(_04826_),
    .A2(_05600_),
    .B1(_05608_),
    .Y(_00540_));
 sky130_fd_sc_hd__nand2_1 _16328_ (.A(net131),
    .B(_05600_),
    .Y(_05609_));
 sky130_fd_sc_hd__o21ai_0 _16329_ (.A1(_04834_),
    .A2(_05600_),
    .B1(_05609_),
    .Y(_00541_));
 sky130_fd_sc_hd__nand2_1 _16330_ (.A(net130),
    .B(_05600_),
    .Y(_05610_));
 sky130_fd_sc_hd__o21ai_0 _16331_ (.A1(_04843_),
    .A2(_05600_),
    .B1(_05610_),
    .Y(_00542_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1271 ();
 sky130_fd_sc_hd__nand2_1 _16333_ (.A(net129),
    .B(_05600_),
    .Y(_05612_));
 sky130_fd_sc_hd__o21ai_0 _16334_ (.A1(_04852_),
    .A2(_05600_),
    .B1(_05612_),
    .Y(_00543_));
 sky130_fd_sc_hd__nand2_1 _16335_ (.A(net128),
    .B(_05600_),
    .Y(_05613_));
 sky130_fd_sc_hd__o21ai_0 _16336_ (.A1(_04860_),
    .A2(_05600_),
    .B1(_05613_),
    .Y(_00544_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1270 ();
 sky130_fd_sc_hd__nand2_1 _16338_ (.A(net127),
    .B(_05600_),
    .Y(_05615_));
 sky130_fd_sc_hd__o21ai_0 _16339_ (.A1(_04871_),
    .A2(_05600_),
    .B1(_05615_),
    .Y(_00514_));
 sky130_fd_sc_hd__nand2_1 _16340_ (.A(net126),
    .B(_05600_),
    .Y(_05616_));
 sky130_fd_sc_hd__o21ai_0 _16341_ (.A1(_04883_),
    .A2(_05600_),
    .B1(_05616_),
    .Y(_00515_));
 sky130_fd_sc_hd__nand2_1 _16342_ (.A(net125),
    .B(_05600_),
    .Y(_05617_));
 sky130_fd_sc_hd__o21ai_0 _16343_ (.A1(_04892_),
    .A2(_05600_),
    .B1(_05617_),
    .Y(_00516_));
 sky130_fd_sc_hd__nand2_1 _16344_ (.A(net124),
    .B(_05600_),
    .Y(_05618_));
 sky130_fd_sc_hd__o21ai_0 _16345_ (.A1(_04899_),
    .A2(_05600_),
    .B1(_05618_),
    .Y(_00517_));
 sky130_fd_sc_hd__nand2_1 _16346_ (.A(net122),
    .B(_05600_),
    .Y(_05619_));
 sky130_fd_sc_hd__o21ai_0 _16347_ (.A1(_04906_),
    .A2(_05600_),
    .B1(_05619_),
    .Y(_00518_));
 sky130_fd_sc_hd__nand2_1 _16348_ (.A(net121),
    .B(_05600_),
    .Y(_05620_));
 sky130_fd_sc_hd__o21ai_0 _16349_ (.A1(_04913_),
    .A2(_05600_),
    .B1(_05620_),
    .Y(_00519_));
 sky130_fd_sc_hd__nand2_1 _16350_ (.A(net120),
    .B(_05600_),
    .Y(_05621_));
 sky130_fd_sc_hd__o21ai_0 _16351_ (.A1(_04923_),
    .A2(_05600_),
    .B1(_05621_),
    .Y(_00520_));
 sky130_fd_sc_hd__nand2_1 _16352_ (.A(net119),
    .B(_05600_),
    .Y(_05622_));
 sky130_fd_sc_hd__o21ai_0 _16353_ (.A1(_04932_),
    .A2(_05600_),
    .B1(_05622_),
    .Y(_00521_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1269 ();
 sky130_fd_sc_hd__nand2_1 _16355_ (.A(net118),
    .B(_05600_),
    .Y(_05624_));
 sky130_fd_sc_hd__o21ai_0 _16356_ (.A1(_04939_),
    .A2(_05600_),
    .B1(_05624_),
    .Y(_00522_));
 sky130_fd_sc_hd__nand2_1 _16357_ (.A(net117),
    .B(_05600_),
    .Y(_05625_));
 sky130_fd_sc_hd__o21ai_0 _16358_ (.A1(_04951_),
    .A2(_05600_),
    .B1(_05625_),
    .Y(_00523_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1268 ();
 sky130_fd_sc_hd__nand2_1 _16360_ (.A(net116),
    .B(_05600_),
    .Y(_05627_));
 sky130_fd_sc_hd__o21ai_0 _16361_ (.A1(_04960_),
    .A2(_05600_),
    .B1(_05627_),
    .Y(_00525_));
 sky130_fd_sc_hd__nand2_1 _16362_ (.A(net115),
    .B(_05600_),
    .Y(_05628_));
 sky130_fd_sc_hd__o21ai_0 _16363_ (.A1(_04974_),
    .A2(_05600_),
    .B1(_05628_),
    .Y(_00526_));
 sky130_fd_sc_hd__nand2_1 _16364_ (.A(net114),
    .B(_05600_),
    .Y(_05629_));
 sky130_fd_sc_hd__o21ai_0 _16365_ (.A1(_04984_),
    .A2(_05600_),
    .B1(_05629_),
    .Y(_00527_));
 sky130_fd_sc_hd__nand2_1 _16366_ (.A(net113),
    .B(_05600_),
    .Y(_05630_));
 sky130_fd_sc_hd__o21ai_0 _16367_ (.A1(_04990_),
    .A2(_05600_),
    .B1(_05630_),
    .Y(_00528_));
 sky130_fd_sc_hd__nand2_1 _16368_ (.A(net110),
    .B(_05600_),
    .Y(_05631_));
 sky130_fd_sc_hd__o21ai_0 _16369_ (.A1(net1129),
    .A2(_05600_),
    .B1(_05631_),
    .Y(_00529_));
 sky130_fd_sc_hd__nand2_1 _16370_ (.A(net109),
    .B(_05600_),
    .Y(_05632_));
 sky130_fd_sc_hd__o21ai_0 _16371_ (.A1(_05011_),
    .A2(_05600_),
    .B1(_05632_),
    .Y(_00530_));
 sky130_fd_sc_hd__nand2_1 _16372_ (.A(net108),
    .B(_05600_),
    .Y(_05633_));
 sky130_fd_sc_hd__o21ai_0 _16373_ (.A1(_05020_),
    .A2(_05600_),
    .B1(_05633_),
    .Y(_00531_));
 sky130_fd_sc_hd__nand2_1 _16374_ (.A(net107),
    .B(_05600_),
    .Y(_05634_));
 sky130_fd_sc_hd__o21ai_0 _16375_ (.A1(_05029_),
    .A2(_05600_),
    .B1(_05634_),
    .Y(_00532_));
 sky130_fd_sc_hd__nand2_1 _16376_ (.A(net106),
    .B(_05600_),
    .Y(_05635_));
 sky130_fd_sc_hd__o21ai_0 _16377_ (.A1(_05035_),
    .A2(_05600_),
    .B1(_05635_),
    .Y(_00533_));
 sky130_fd_sc_hd__nand2_1 _16378_ (.A(net105),
    .B(_05600_),
    .Y(_05636_));
 sky130_fd_sc_hd__o21ai_0 _16379_ (.A1(_05044_),
    .A2(_05600_),
    .B1(_05636_),
    .Y(_00534_));
 sky130_fd_sc_hd__nand2_1 _16380_ (.A(net104),
    .B(_05600_),
    .Y(_05637_));
 sky130_fd_sc_hd__o21ai_0 _16381_ (.A1(_05060_),
    .A2(_05600_),
    .B1(_05637_),
    .Y(_00536_));
 sky130_fd_sc_hd__mux2i_1 _16382_ (.A0(_05113_),
    .A1(net103),
    .S(_05600_),
    .Y(_05638_));
 sky130_fd_sc_hd__o21ai_0 _16383_ (.A1(_05112_),
    .A2(_05600_),
    .B1(_05638_),
    .Y(_00537_));
 sky130_fd_sc_hd__nor4_4 _16384_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(net1039),
    .D(_09803_),
    .Y(_05639_));
 sky130_fd_sc_hd__nor2_1 _16385_ (.A(net173),
    .B(_05639_),
    .Y(_05640_));
 sky130_fd_sc_hd__a21oi_1 _16386_ (.A1(_05118_),
    .A2(_05639_),
    .B1(_05640_),
    .Y(_00545_));
 sky130_fd_sc_hd__nor2_1 _16387_ (.A(net172),
    .B(_05639_),
    .Y(_05641_));
 sky130_fd_sc_hd__a21oi_1 _16388_ (.A1(_05122_),
    .A2(_05639_),
    .B1(_05641_),
    .Y(_00556_));
 sky130_fd_sc_hd__nand2_8 _16389_ (.A(_09731_),
    .B(_09836_),
    .Y(_05642_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1266 ();
 sky130_fd_sc_hd__nand2_1 _16392_ (.A(net171),
    .B(_05642_),
    .Y(_05645_));
 sky130_fd_sc_hd__o21ai_0 _16393_ (.A1(_05126_),
    .A2(_05642_),
    .B1(_05645_),
    .Y(_00567_));
 sky130_fd_sc_hd__nor2_1 _16394_ (.A(net170),
    .B(_05639_),
    .Y(_05646_));
 sky130_fd_sc_hd__a21oi_1 _16395_ (.A1(_05132_),
    .A2(_05639_),
    .B1(_05646_),
    .Y(_00570_));
 sky130_fd_sc_hd__nand2_1 _16396_ (.A(net169),
    .B(_05642_),
    .Y(_05647_));
 sky130_fd_sc_hd__o21ai_0 _16397_ (.A1(_05140_),
    .A2(_05642_),
    .B1(_05647_),
    .Y(_00571_));
 sky130_fd_sc_hd__nand2_1 _16398_ (.A(net168),
    .B(_05642_),
    .Y(_05648_));
 sky130_fd_sc_hd__o21ai_0 _16399_ (.A1(_05149_),
    .A2(_05642_),
    .B1(_05648_),
    .Y(_00572_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1265 ();
 sky130_fd_sc_hd__nand2_1 _16401_ (.A(net166),
    .B(_05642_),
    .Y(_05650_));
 sky130_fd_sc_hd__o21ai_0 _16402_ (.A1(_05157_),
    .A2(_05642_),
    .B1(_05650_),
    .Y(_00573_));
 sky130_fd_sc_hd__nand2_1 _16403_ (.A(net165),
    .B(_05642_),
    .Y(_05651_));
 sky130_fd_sc_hd__o21ai_0 _16404_ (.A1(_05166_),
    .A2(_05642_),
    .B1(_05651_),
    .Y(_00574_));
 sky130_fd_sc_hd__nand2_1 _16405_ (.A(net164),
    .B(_05642_),
    .Y(_05652_));
 sky130_fd_sc_hd__o21ai_0 _16406_ (.A1(_05173_),
    .A2(_05642_),
    .B1(_05652_),
    .Y(_00575_));
 sky130_fd_sc_hd__nand2_1 _16407_ (.A(net163),
    .B(_05642_),
    .Y(_05653_));
 sky130_fd_sc_hd__o21ai_0 _16408_ (.A1(_05183_),
    .A2(_05642_),
    .B1(_05653_),
    .Y(_00576_));
 sky130_fd_sc_hd__nand2_1 _16409_ (.A(net162),
    .B(_05642_),
    .Y(_05654_));
 sky130_fd_sc_hd__o21ai_0 _16410_ (.A1(_05192_),
    .A2(_05642_),
    .B1(_05654_),
    .Y(_00546_));
 sky130_fd_sc_hd__nand2_1 _16411_ (.A(net161),
    .B(_05642_),
    .Y(_05655_));
 sky130_fd_sc_hd__o21ai_0 _16412_ (.A1(_05204_),
    .A2(_05642_),
    .B1(_05655_),
    .Y(_00547_));
 sky130_fd_sc_hd__nand2_1 _16413_ (.A(net160),
    .B(_05642_),
    .Y(_05656_));
 sky130_fd_sc_hd__o21ai_0 _16414_ (.A1(_05214_),
    .A2(_05642_),
    .B1(_05656_),
    .Y(_00548_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1264 ();
 sky130_fd_sc_hd__nand2_1 _16416_ (.A(net159),
    .B(_05642_),
    .Y(_05658_));
 sky130_fd_sc_hd__o21ai_0 _16417_ (.A1(_05221_),
    .A2(_05642_),
    .B1(_05658_),
    .Y(_00549_));
 sky130_fd_sc_hd__nand2_1 _16418_ (.A(net158),
    .B(_05642_),
    .Y(_05659_));
 sky130_fd_sc_hd__o21ai_0 _16419_ (.A1(_05228_),
    .A2(_05642_),
    .B1(_05659_),
    .Y(_00550_));
 sky130_fd_sc_hd__nand2_1 _16420_ (.A(net157),
    .B(_05642_),
    .Y(_05660_));
 sky130_fd_sc_hd__o21ai_0 _16421_ (.A1(_05238_),
    .A2(_05642_),
    .B1(_05660_),
    .Y(_00551_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1263 ();
 sky130_fd_sc_hd__nand2_1 _16423_ (.A(net155),
    .B(_05642_),
    .Y(_05662_));
 sky130_fd_sc_hd__o21ai_0 _16424_ (.A1(_05247_),
    .A2(_05642_),
    .B1(_05662_),
    .Y(_00552_));
 sky130_fd_sc_hd__nand2_1 _16425_ (.A(net154),
    .B(_05642_),
    .Y(_05663_));
 sky130_fd_sc_hd__o21ai_0 _16426_ (.A1(_05258_),
    .A2(_05642_),
    .B1(_05663_),
    .Y(_00553_));
 sky130_fd_sc_hd__nand2_1 _16427_ (.A(net153),
    .B(_05642_),
    .Y(_05664_));
 sky130_fd_sc_hd__o21ai_0 _16428_ (.A1(_05267_),
    .A2(_05642_),
    .B1(_05664_),
    .Y(_00554_));
 sky130_fd_sc_hd__nand2_1 _16429_ (.A(net152),
    .B(_05642_),
    .Y(_05665_));
 sky130_fd_sc_hd__o21ai_0 _16430_ (.A1(_05280_),
    .A2(_05642_),
    .B1(_05665_),
    .Y(_00555_));
 sky130_fd_sc_hd__nand2_1 _16431_ (.A(net151),
    .B(_05642_),
    .Y(_05666_));
 sky130_fd_sc_hd__o21ai_0 _16432_ (.A1(_05291_),
    .A2(_05642_),
    .B1(_05666_),
    .Y(_00557_));
 sky130_fd_sc_hd__nand2_1 _16433_ (.A(net150),
    .B(_05642_),
    .Y(_05667_));
 sky130_fd_sc_hd__o21ai_0 _16434_ (.A1(_05301_),
    .A2(_05642_),
    .B1(_05667_),
    .Y(_00558_));
 sky130_fd_sc_hd__nand2_1 _16435_ (.A(net149),
    .B(_05642_),
    .Y(_05668_));
 sky130_fd_sc_hd__o21ai_0 _16436_ (.A1(_05309_),
    .A2(_05642_),
    .B1(_05668_),
    .Y(_00559_));
 sky130_fd_sc_hd__nand2_1 _16437_ (.A(net148),
    .B(_05642_),
    .Y(_05669_));
 sky130_fd_sc_hd__o21ai_0 _16438_ (.A1(_05320_),
    .A2(_05642_),
    .B1(_05669_),
    .Y(_00560_));
 sky130_fd_sc_hd__nand2_1 _16439_ (.A(net147),
    .B(_05642_),
    .Y(_05670_));
 sky130_fd_sc_hd__o21ai_0 _16440_ (.A1(net1145),
    .A2(_05642_),
    .B1(_05670_),
    .Y(_00561_));
 sky130_fd_sc_hd__nand2_1 _16441_ (.A(net146),
    .B(_05642_),
    .Y(_05671_));
 sky130_fd_sc_hd__o21ai_0 _16442_ (.A1(_05339_),
    .A2(_05642_),
    .B1(_05671_),
    .Y(_00562_));
 sky130_fd_sc_hd__nand2_1 _16443_ (.A(net144),
    .B(_05642_),
    .Y(_05672_));
 sky130_fd_sc_hd__o21ai_0 _16444_ (.A1(_05347_),
    .A2(_05642_),
    .B1(_05672_),
    .Y(_00563_));
 sky130_fd_sc_hd__nor2_1 _16445_ (.A(net143),
    .B(_05639_),
    .Y(_05673_));
 sky130_fd_sc_hd__a21oi_1 _16446_ (.A1(_05358_),
    .A2(_05639_),
    .B1(_05673_),
    .Y(_00564_));
 sky130_fd_sc_hd__nand2_1 _16447_ (.A(net142),
    .B(_05642_),
    .Y(_05674_));
 sky130_fd_sc_hd__o21ai_0 _16448_ (.A1(_05372_),
    .A2(_05642_),
    .B1(_05674_),
    .Y(_00565_));
 sky130_fd_sc_hd__nand2_1 _16449_ (.A(net141),
    .B(_05642_),
    .Y(_05675_));
 sky130_fd_sc_hd__o21ai_0 _16450_ (.A1(_05380_),
    .A2(_05642_),
    .B1(_05675_),
    .Y(_00566_));
 sky130_fd_sc_hd__nor2_1 _16451_ (.A(net140),
    .B(_05639_),
    .Y(_05676_));
 sky130_fd_sc_hd__a21oi_1 _16452_ (.A1(net1143),
    .A2(_05639_),
    .B1(_05676_),
    .Y(_00568_));
 sky130_fd_sc_hd__nand2_1 _16453_ (.A(net139),
    .B(_05642_),
    .Y(_05677_));
 sky130_fd_sc_hd__o21ai_0 _16454_ (.A1(_05430_),
    .A2(_05642_),
    .B1(_05677_),
    .Y(_00569_));
 sky130_fd_sc_hd__nand2_8 _16455_ (.A(_09739_),
    .B(_04784_),
    .Y(_05678_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1261 ();
 sky130_fd_sc_hd__nand2_1 _16458_ (.A(net208),
    .B(_05678_),
    .Y(_05681_));
 sky130_fd_sc_hd__o21ai_0 _16459_ (.A1(_04790_),
    .A2(_05678_),
    .B1(_05681_),
    .Y(_00577_));
 sky130_fd_sc_hd__nand2_1 _16460_ (.A(net207),
    .B(_05678_),
    .Y(_05682_));
 sky130_fd_sc_hd__o21ai_0 _16461_ (.A1(_04794_),
    .A2(_05678_),
    .B1(_05682_),
    .Y(_00588_));
 sky130_fd_sc_hd__nand2_1 _16462_ (.A(net206),
    .B(_05678_),
    .Y(_05683_));
 sky130_fd_sc_hd__o21ai_0 _16463_ (.A1(_04801_),
    .A2(_05678_),
    .B1(_05683_),
    .Y(_00599_));
 sky130_fd_sc_hd__nand2_1 _16464_ (.A(net205),
    .B(_05678_),
    .Y(_05684_));
 sky130_fd_sc_hd__o21ai_0 _16465_ (.A1(_04808_),
    .A2(_05678_),
    .B1(_05684_),
    .Y(_00602_));
 sky130_fd_sc_hd__nand2_1 _16466_ (.A(net204),
    .B(_05678_),
    .Y(_05685_));
 sky130_fd_sc_hd__o21ai_0 _16467_ (.A1(_04817_),
    .A2(_05678_),
    .B1(_05685_),
    .Y(_00603_));
 sky130_fd_sc_hd__nand2_1 _16468_ (.A(net203),
    .B(_05678_),
    .Y(_05686_));
 sky130_fd_sc_hd__o21ai_0 _16469_ (.A1(_04826_),
    .A2(_05678_),
    .B1(_05686_),
    .Y(_00604_));
 sky130_fd_sc_hd__nand2_1 _16470_ (.A(net202),
    .B(_05678_),
    .Y(_05687_));
 sky130_fd_sc_hd__o21ai_0 _16471_ (.A1(_04834_),
    .A2(_05678_),
    .B1(_05687_),
    .Y(_00605_));
 sky130_fd_sc_hd__nand2_1 _16472_ (.A(net201),
    .B(_05678_),
    .Y(_05688_));
 sky130_fd_sc_hd__o21ai_0 _16473_ (.A1(_04843_),
    .A2(_05678_),
    .B1(_05688_),
    .Y(_00606_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1260 ();
 sky130_fd_sc_hd__nand2_1 _16475_ (.A(net199),
    .B(_05678_),
    .Y(_05690_));
 sky130_fd_sc_hd__o21ai_0 _16476_ (.A1(_04852_),
    .A2(_05678_),
    .B1(_05690_),
    .Y(_00607_));
 sky130_fd_sc_hd__nand2_1 _16477_ (.A(net198),
    .B(_05678_),
    .Y(_05691_));
 sky130_fd_sc_hd__o21ai_0 _16478_ (.A1(_04860_),
    .A2(_05678_),
    .B1(_05691_),
    .Y(_00608_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1259 ();
 sky130_fd_sc_hd__nand2_1 _16480_ (.A(net197),
    .B(_05678_),
    .Y(_05693_));
 sky130_fd_sc_hd__o21ai_0 _16481_ (.A1(_04871_),
    .A2(_05678_),
    .B1(_05693_),
    .Y(_00578_));
 sky130_fd_sc_hd__nand2_1 _16482_ (.A(net196),
    .B(_05678_),
    .Y(_05694_));
 sky130_fd_sc_hd__o21ai_0 _16483_ (.A1(_04883_),
    .A2(_05678_),
    .B1(_05694_),
    .Y(_00579_));
 sky130_fd_sc_hd__nand2_1 _16484_ (.A(net195),
    .B(_05678_),
    .Y(_05695_));
 sky130_fd_sc_hd__o21ai_0 _16485_ (.A1(_04892_),
    .A2(_05678_),
    .B1(_05695_),
    .Y(_00580_));
 sky130_fd_sc_hd__nand2_1 _16486_ (.A(net194),
    .B(_05678_),
    .Y(_05696_));
 sky130_fd_sc_hd__o21ai_0 _16487_ (.A1(_04899_),
    .A2(_05678_),
    .B1(_05696_),
    .Y(_00581_));
 sky130_fd_sc_hd__nand2_1 _16488_ (.A(net193),
    .B(_05678_),
    .Y(_05697_));
 sky130_fd_sc_hd__o21ai_0 _16489_ (.A1(_04906_),
    .A2(_05678_),
    .B1(_05697_),
    .Y(_00582_));
 sky130_fd_sc_hd__nand2_1 _16490_ (.A(net192),
    .B(_05678_),
    .Y(_05698_));
 sky130_fd_sc_hd__o21ai_0 _16491_ (.A1(_04913_),
    .A2(_05678_),
    .B1(_05698_),
    .Y(_00583_));
 sky130_fd_sc_hd__nand2_1 _16492_ (.A(net191),
    .B(_05678_),
    .Y(_05699_));
 sky130_fd_sc_hd__o21ai_0 _16493_ (.A1(_04923_),
    .A2(_05678_),
    .B1(_05699_),
    .Y(_00584_));
 sky130_fd_sc_hd__nand2_1 _16494_ (.A(net190),
    .B(_05678_),
    .Y(_05700_));
 sky130_fd_sc_hd__o21ai_0 _16495_ (.A1(_04932_),
    .A2(_05678_),
    .B1(_05700_),
    .Y(_00585_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1258 ();
 sky130_fd_sc_hd__nand2_1 _16497_ (.A(net188),
    .B(_05678_),
    .Y(_05702_));
 sky130_fd_sc_hd__o21ai_0 _16498_ (.A1(_04939_),
    .A2(_05678_),
    .B1(_05702_),
    .Y(_00586_));
 sky130_fd_sc_hd__nand2_1 _16499_ (.A(net187),
    .B(_05678_),
    .Y(_05703_));
 sky130_fd_sc_hd__o21ai_0 _16500_ (.A1(_04951_),
    .A2(_05678_),
    .B1(_05703_),
    .Y(_00587_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1257 ();
 sky130_fd_sc_hd__nand2_1 _16502_ (.A(net186),
    .B(_05678_),
    .Y(_05705_));
 sky130_fd_sc_hd__o21ai_0 _16503_ (.A1(_04960_),
    .A2(_05678_),
    .B1(_05705_),
    .Y(_00589_));
 sky130_fd_sc_hd__nand2_1 _16504_ (.A(net185),
    .B(_05678_),
    .Y(_05706_));
 sky130_fd_sc_hd__o21ai_0 _16505_ (.A1(_04974_),
    .A2(_05678_),
    .B1(_05706_),
    .Y(_00590_));
 sky130_fd_sc_hd__nand2_1 _16506_ (.A(net184),
    .B(_05678_),
    .Y(_05707_));
 sky130_fd_sc_hd__o21ai_0 _16507_ (.A1(_04984_),
    .A2(_05678_),
    .B1(_05707_),
    .Y(_00591_));
 sky130_fd_sc_hd__nand2_1 _16508_ (.A(net183),
    .B(_05678_),
    .Y(_05708_));
 sky130_fd_sc_hd__o21ai_0 _16509_ (.A1(_04990_),
    .A2(_05678_),
    .B1(_05708_),
    .Y(_00592_));
 sky130_fd_sc_hd__nand2_1 _16510_ (.A(net182),
    .B(_05678_),
    .Y(_05709_));
 sky130_fd_sc_hd__o21ai_0 _16511_ (.A1(net1129),
    .A2(_05678_),
    .B1(_05709_),
    .Y(_00593_));
 sky130_fd_sc_hd__nand2_1 _16512_ (.A(net181),
    .B(_05678_),
    .Y(_05710_));
 sky130_fd_sc_hd__o21ai_0 _16513_ (.A1(_05011_),
    .A2(_05678_),
    .B1(_05710_),
    .Y(_00594_));
 sky130_fd_sc_hd__nand2_1 _16514_ (.A(net180),
    .B(_05678_),
    .Y(_05711_));
 sky130_fd_sc_hd__o21ai_0 _16515_ (.A1(_05020_),
    .A2(_05678_),
    .B1(_05711_),
    .Y(_00595_));
 sky130_fd_sc_hd__nand2_1 _16516_ (.A(net179),
    .B(_05678_),
    .Y(_05712_));
 sky130_fd_sc_hd__o21ai_0 _16517_ (.A1(_05029_),
    .A2(_05678_),
    .B1(_05712_),
    .Y(_00596_));
 sky130_fd_sc_hd__nand2_1 _16518_ (.A(net177),
    .B(_05678_),
    .Y(_05713_));
 sky130_fd_sc_hd__o21ai_0 _16519_ (.A1(_05035_),
    .A2(_05678_),
    .B1(_05713_),
    .Y(_00597_));
 sky130_fd_sc_hd__nand2_1 _16520_ (.A(net176),
    .B(_05678_),
    .Y(_05714_));
 sky130_fd_sc_hd__o21ai_0 _16521_ (.A1(_05044_),
    .A2(_05678_),
    .B1(_05714_),
    .Y(_00598_));
 sky130_fd_sc_hd__nand2_1 _16522_ (.A(net175),
    .B(_05678_),
    .Y(_05715_));
 sky130_fd_sc_hd__o21ai_0 _16523_ (.A1(_05060_),
    .A2(_05678_),
    .B1(_05715_),
    .Y(_00600_));
 sky130_fd_sc_hd__mux2i_1 _16524_ (.A0(_05113_),
    .A1(net174),
    .S(_05678_),
    .Y(_05716_));
 sky130_fd_sc_hd__o21ai_0 _16525_ (.A1(_05112_),
    .A2(_05678_),
    .B1(_05716_),
    .Y(_00601_));
 sky130_fd_sc_hd__nand2_8 _16526_ (.A(net551),
    .B(_05115_),
    .Y(_05717_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1255 ();
 sky130_fd_sc_hd__nand2_1 _16529_ (.A(net244),
    .B(_05717_),
    .Y(_05720_));
 sky130_fd_sc_hd__o21ai_0 _16530_ (.A1(_05118_),
    .A2(_05717_),
    .B1(_05720_),
    .Y(_00609_));
 sky130_fd_sc_hd__nand2_1 _16531_ (.A(net243),
    .B(_05717_),
    .Y(_05721_));
 sky130_fd_sc_hd__o21ai_0 _16532_ (.A1(_05122_),
    .A2(_05717_),
    .B1(_05721_),
    .Y(_00620_));
 sky130_fd_sc_hd__nand2_1 _16533_ (.A(net242),
    .B(_05717_),
    .Y(_05722_));
 sky130_fd_sc_hd__o21ai_0 _16534_ (.A1(_05126_),
    .A2(_05717_),
    .B1(_05722_),
    .Y(_00631_));
 sky130_fd_sc_hd__nand2_1 _16535_ (.A(net241),
    .B(_05717_),
    .Y(_05723_));
 sky130_fd_sc_hd__o21ai_0 _16536_ (.A1(_05132_),
    .A2(_05717_),
    .B1(_05723_),
    .Y(_00634_));
 sky130_fd_sc_hd__nand2_1 _16537_ (.A(net240),
    .B(_05717_),
    .Y(_05724_));
 sky130_fd_sc_hd__o21ai_0 _16538_ (.A1(_05140_),
    .A2(_05717_),
    .B1(_05724_),
    .Y(_00635_));
 sky130_fd_sc_hd__nand2_1 _16539_ (.A(net239),
    .B(_05717_),
    .Y(_05725_));
 sky130_fd_sc_hd__o21ai_0 _16540_ (.A1(_05149_),
    .A2(_05717_),
    .B1(_05725_),
    .Y(_00636_));
 sky130_fd_sc_hd__nand2_1 _16541_ (.A(net238),
    .B(_05717_),
    .Y(_05726_));
 sky130_fd_sc_hd__o21ai_0 _16542_ (.A1(_05157_),
    .A2(_05717_),
    .B1(_05726_),
    .Y(_00637_));
 sky130_fd_sc_hd__nand2_1 _16543_ (.A(net237),
    .B(_05717_),
    .Y(_05727_));
 sky130_fd_sc_hd__o21ai_0 _16544_ (.A1(_05166_),
    .A2(_05717_),
    .B1(_05727_),
    .Y(_00638_));
 sky130_fd_sc_hd__nand2_1 _16545_ (.A(net236),
    .B(_05717_),
    .Y(_05728_));
 sky130_fd_sc_hd__o21ai_0 _16546_ (.A1(_05173_),
    .A2(_05717_),
    .B1(_05728_),
    .Y(_00639_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1254 ();
 sky130_fd_sc_hd__nand2_2 _16548_ (.A(net235),
    .B(_05717_),
    .Y(_05730_));
 sky130_fd_sc_hd__o21ai_0 _16549_ (.A1(_05183_),
    .A2(_05717_),
    .B1(_05730_),
    .Y(_00640_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1253 ();
 sky130_fd_sc_hd__nand2_1 _16551_ (.A(net233),
    .B(_05717_),
    .Y(_05732_));
 sky130_fd_sc_hd__o21ai_0 _16552_ (.A1(_05192_),
    .A2(_05717_),
    .B1(_05732_),
    .Y(_00610_));
 sky130_fd_sc_hd__nand2_1 _16553_ (.A(net232),
    .B(_05717_),
    .Y(_05733_));
 sky130_fd_sc_hd__o21ai_0 _16554_ (.A1(_05204_),
    .A2(_05717_),
    .B1(_05733_),
    .Y(_00611_));
 sky130_fd_sc_hd__nand2_1 _16555_ (.A(net231),
    .B(_05717_),
    .Y(_05734_));
 sky130_fd_sc_hd__o21ai_0 _16556_ (.A1(_05214_),
    .A2(_05717_),
    .B1(_05734_),
    .Y(_00612_));
 sky130_fd_sc_hd__nand2_1 _16557_ (.A(net230),
    .B(_05717_),
    .Y(_05735_));
 sky130_fd_sc_hd__o21ai_0 _16558_ (.A1(_05221_),
    .A2(_05717_),
    .B1(_05735_),
    .Y(_00613_));
 sky130_fd_sc_hd__nand2_1 _16559_ (.A(net229),
    .B(_05717_),
    .Y(_05736_));
 sky130_fd_sc_hd__o21ai_0 _16560_ (.A1(_05228_),
    .A2(_05717_),
    .B1(_05736_),
    .Y(_00614_));
 sky130_fd_sc_hd__nand2_1 _16561_ (.A(net228),
    .B(_05717_),
    .Y(_05737_));
 sky130_fd_sc_hd__o21ai_0 _16562_ (.A1(_05238_),
    .A2(_05717_),
    .B1(_05737_),
    .Y(_00615_));
 sky130_fd_sc_hd__nand2_1 _16563_ (.A(net227),
    .B(_05717_),
    .Y(_05738_));
 sky130_fd_sc_hd__o21ai_0 _16564_ (.A1(_05247_),
    .A2(_05717_),
    .B1(_05738_),
    .Y(_00616_));
 sky130_fd_sc_hd__nand2_1 _16565_ (.A(net226),
    .B(_05717_),
    .Y(_05739_));
 sky130_fd_sc_hd__o21ai_0 _16566_ (.A1(_05258_),
    .A2(_05717_),
    .B1(_05739_),
    .Y(_00617_));
 sky130_fd_sc_hd__nand2_1 _16567_ (.A(net225),
    .B(_05717_),
    .Y(_05740_));
 sky130_fd_sc_hd__o21ai_0 _16568_ (.A1(_05267_),
    .A2(_05717_),
    .B1(_05740_),
    .Y(_00618_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1252 ();
 sky130_fd_sc_hd__nand2_1 _16570_ (.A(net224),
    .B(_05717_),
    .Y(_05742_));
 sky130_fd_sc_hd__o21ai_0 _16571_ (.A1(_05280_),
    .A2(_05717_),
    .B1(_05742_),
    .Y(_00619_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1251 ();
 sky130_fd_sc_hd__nand2_1 _16573_ (.A(net221),
    .B(_05717_),
    .Y(_05744_));
 sky130_fd_sc_hd__o21ai_0 _16574_ (.A1(_05291_),
    .A2(_05717_),
    .B1(_05744_),
    .Y(_00621_));
 sky130_fd_sc_hd__nand2_1 _16575_ (.A(net220),
    .B(_05717_),
    .Y(_05745_));
 sky130_fd_sc_hd__o21ai_0 _16576_ (.A1(_05301_),
    .A2(_05717_),
    .B1(_05745_),
    .Y(_00622_));
 sky130_fd_sc_hd__nand2_1 _16577_ (.A(net219),
    .B(_05717_),
    .Y(_05746_));
 sky130_fd_sc_hd__o21ai_0 _16578_ (.A1(_05309_),
    .A2(_05717_),
    .B1(_05746_),
    .Y(_00623_));
 sky130_fd_sc_hd__nand2_1 _16579_ (.A(net218),
    .B(_05717_),
    .Y(_05747_));
 sky130_fd_sc_hd__o21ai_0 _16580_ (.A1(_05320_),
    .A2(_05717_),
    .B1(_05747_),
    .Y(_00624_));
 sky130_fd_sc_hd__nand2_1 _16581_ (.A(net217),
    .B(_05717_),
    .Y(_05748_));
 sky130_fd_sc_hd__o21ai_0 _16582_ (.A1(net1145),
    .A2(_05717_),
    .B1(_05748_),
    .Y(_00625_));
 sky130_fd_sc_hd__nand2_1 _16583_ (.A(net216),
    .B(_05717_),
    .Y(_05749_));
 sky130_fd_sc_hd__o21ai_0 _16584_ (.A1(_05339_),
    .A2(_05717_),
    .B1(_05749_),
    .Y(_00626_));
 sky130_fd_sc_hd__nand2_1 _16585_ (.A(net215),
    .B(_05717_),
    .Y(_05750_));
 sky130_fd_sc_hd__o21ai_0 _16586_ (.A1(_05347_),
    .A2(_05717_),
    .B1(_05750_),
    .Y(_00627_));
 sky130_fd_sc_hd__nand2_1 _16587_ (.A(net214),
    .B(_05717_),
    .Y(_05751_));
 sky130_fd_sc_hd__o21ai_0 _16588_ (.A1(_05358_),
    .A2(_05717_),
    .B1(_05751_),
    .Y(_00628_));
 sky130_fd_sc_hd__nand2_1 _16589_ (.A(net213),
    .B(_05717_),
    .Y(_05752_));
 sky130_fd_sc_hd__o21ai_0 _16590_ (.A1(_05372_),
    .A2(_05717_),
    .B1(_05752_),
    .Y(_00629_));
 sky130_fd_sc_hd__nand2_1 _16591_ (.A(net212),
    .B(_05717_),
    .Y(_05753_));
 sky130_fd_sc_hd__o21ai_0 _16592_ (.A1(_05380_),
    .A2(_05717_),
    .B1(_05753_),
    .Y(_00630_));
 sky130_fd_sc_hd__a21oi_1 _16593_ (.A1(_09784_),
    .A2(_05115_),
    .B1(net210),
    .Y(_05754_));
 sky130_fd_sc_hd__a31oi_1 _16594_ (.A1(_09784_),
    .A2(_05115_),
    .A3(net1143),
    .B1(_05754_),
    .Y(_00632_));
 sky130_fd_sc_hd__nand2_1 _16595_ (.A(net209),
    .B(_05717_),
    .Y(_05755_));
 sky130_fd_sc_hd__o21ai_0 _16596_ (.A1(_05430_),
    .A2(_05717_),
    .B1(_05755_),
    .Y(_00633_));
 sky130_fd_sc_hd__nand2_8 _16597_ (.A(_09739_),
    .B(_05433_),
    .Y(_05756_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1249 ();
 sky130_fd_sc_hd__nand2_1 _16600_ (.A(net280),
    .B(_05756_),
    .Y(_05759_));
 sky130_fd_sc_hd__o21ai_0 _16601_ (.A1(_04790_),
    .A2(_05756_),
    .B1(_05759_),
    .Y(_00161_));
 sky130_fd_sc_hd__nand2_1 _16602_ (.A(net279),
    .B(_05756_),
    .Y(_05760_));
 sky130_fd_sc_hd__o21ai_0 _16603_ (.A1(_04794_),
    .A2(_05756_),
    .B1(_05760_),
    .Y(_00172_));
 sky130_fd_sc_hd__nand2_1 _16604_ (.A(net277),
    .B(_05756_),
    .Y(_05761_));
 sky130_fd_sc_hd__o21ai_0 _16605_ (.A1(_04801_),
    .A2(_05756_),
    .B1(_05761_),
    .Y(_00183_));
 sky130_fd_sc_hd__nand2_1 _16606_ (.A(net276),
    .B(_05756_),
    .Y(_05762_));
 sky130_fd_sc_hd__o21ai_0 _16607_ (.A1(_04808_),
    .A2(_05756_),
    .B1(_05762_),
    .Y(_00186_));
 sky130_fd_sc_hd__nand2_1 _16608_ (.A(net275),
    .B(_05756_),
    .Y(_05763_));
 sky130_fd_sc_hd__o21ai_0 _16609_ (.A1(_04817_),
    .A2(_05756_),
    .B1(_05763_),
    .Y(_00187_));
 sky130_fd_sc_hd__nand2_1 _16610_ (.A(net274),
    .B(_05756_),
    .Y(_05764_));
 sky130_fd_sc_hd__o21ai_0 _16611_ (.A1(_04826_),
    .A2(_05756_),
    .B1(_05764_),
    .Y(_00188_));
 sky130_fd_sc_hd__nand2_1 _16612_ (.A(net273),
    .B(_05756_),
    .Y(_05765_));
 sky130_fd_sc_hd__o21ai_0 _16613_ (.A1(_04834_),
    .A2(_05756_),
    .B1(_05765_),
    .Y(_00189_));
 sky130_fd_sc_hd__nand2_1 _16614_ (.A(net272),
    .B(_05756_),
    .Y(_05766_));
 sky130_fd_sc_hd__o21ai_0 _16615_ (.A1(_04843_),
    .A2(_05756_),
    .B1(_05766_),
    .Y(_00190_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1248 ();
 sky130_fd_sc_hd__nand2_1 _16617_ (.A(net271),
    .B(_05756_),
    .Y(_05768_));
 sky130_fd_sc_hd__o21ai_0 _16618_ (.A1(_04852_),
    .A2(_05756_),
    .B1(_05768_),
    .Y(_00191_));
 sky130_fd_sc_hd__nand2_1 _16619_ (.A(net270),
    .B(_05756_),
    .Y(_05769_));
 sky130_fd_sc_hd__o21ai_0 _16620_ (.A1(_04860_),
    .A2(_05756_),
    .B1(_05769_),
    .Y(_00192_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1247 ();
 sky130_fd_sc_hd__nand2_1 _16622_ (.A(net269),
    .B(_05756_),
    .Y(_05771_));
 sky130_fd_sc_hd__o21ai_0 _16623_ (.A1(_04871_),
    .A2(_05756_),
    .B1(_05771_),
    .Y(_00162_));
 sky130_fd_sc_hd__nand2_1 _16624_ (.A(net268),
    .B(_05756_),
    .Y(_05772_));
 sky130_fd_sc_hd__o21ai_0 _16625_ (.A1(_04883_),
    .A2(_05756_),
    .B1(_05772_),
    .Y(_00163_));
 sky130_fd_sc_hd__nand2_1 _16626_ (.A(net266),
    .B(_05756_),
    .Y(_05773_));
 sky130_fd_sc_hd__o21ai_0 _16627_ (.A1(_04892_),
    .A2(_05756_),
    .B1(_05773_),
    .Y(_00164_));
 sky130_fd_sc_hd__nand2_1 _16628_ (.A(net265),
    .B(_05756_),
    .Y(_05774_));
 sky130_fd_sc_hd__o21ai_0 _16629_ (.A1(_04899_),
    .A2(_05756_),
    .B1(_05774_),
    .Y(_00165_));
 sky130_fd_sc_hd__nand2_1 _16630_ (.A(net264),
    .B(_05756_),
    .Y(_05775_));
 sky130_fd_sc_hd__o21ai_0 _16631_ (.A1(_04906_),
    .A2(_05756_),
    .B1(_05775_),
    .Y(_00166_));
 sky130_fd_sc_hd__nand2_1 _16632_ (.A(net263),
    .B(_05756_),
    .Y(_05776_));
 sky130_fd_sc_hd__o21ai_0 _16633_ (.A1(_04913_),
    .A2(_05756_),
    .B1(_05776_),
    .Y(_00167_));
 sky130_fd_sc_hd__nand2_1 _16634_ (.A(net262),
    .B(_05756_),
    .Y(_05777_));
 sky130_fd_sc_hd__o21ai_0 _16635_ (.A1(_04923_),
    .A2(_05756_),
    .B1(_05777_),
    .Y(_00168_));
 sky130_fd_sc_hd__nand2_1 _16636_ (.A(net261),
    .B(_05756_),
    .Y(_05778_));
 sky130_fd_sc_hd__o21ai_0 _16637_ (.A1(_04932_),
    .A2(_05756_),
    .B1(_05778_),
    .Y(_00169_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1246 ();
 sky130_fd_sc_hd__nand2_1 _16639_ (.A(net260),
    .B(_05756_),
    .Y(_05780_));
 sky130_fd_sc_hd__o21ai_0 _16640_ (.A1(_04939_),
    .A2(_05756_),
    .B1(_05780_),
    .Y(_00170_));
 sky130_fd_sc_hd__nand2_1 _16641_ (.A(net259),
    .B(_05756_),
    .Y(_05781_));
 sky130_fd_sc_hd__o21ai_0 _16642_ (.A1(_04951_),
    .A2(_05756_),
    .B1(_05781_),
    .Y(_00171_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1245 ();
 sky130_fd_sc_hd__nand2_1 _16644_ (.A(net258),
    .B(_05756_),
    .Y(_05783_));
 sky130_fd_sc_hd__o21ai_0 _16645_ (.A1(_04960_),
    .A2(_05756_),
    .B1(_05783_),
    .Y(_00173_));
 sky130_fd_sc_hd__nand2_1 _16646_ (.A(net257),
    .B(_05756_),
    .Y(_05784_));
 sky130_fd_sc_hd__o21ai_0 _16647_ (.A1(_04974_),
    .A2(_05756_),
    .B1(_05784_),
    .Y(_00174_));
 sky130_fd_sc_hd__nand2_1 _16648_ (.A(net255),
    .B(_05756_),
    .Y(_05785_));
 sky130_fd_sc_hd__o21ai_0 _16649_ (.A1(_04984_),
    .A2(_05756_),
    .B1(_05785_),
    .Y(_00175_));
 sky130_fd_sc_hd__nand2_1 _16650_ (.A(net254),
    .B(_05756_),
    .Y(_05786_));
 sky130_fd_sc_hd__o21ai_0 _16651_ (.A1(_04990_),
    .A2(_05756_),
    .B1(_05786_),
    .Y(_00176_));
 sky130_fd_sc_hd__nand2_1 _16652_ (.A(net253),
    .B(_05756_),
    .Y(_05787_));
 sky130_fd_sc_hd__o21ai_0 _16653_ (.A1(net1129),
    .A2(_05756_),
    .B1(_05787_),
    .Y(_00177_));
 sky130_fd_sc_hd__nand2_1 _16654_ (.A(net252),
    .B(_05756_),
    .Y(_05788_));
 sky130_fd_sc_hd__o21ai_0 _16655_ (.A1(_05011_),
    .A2(_05756_),
    .B1(_05788_),
    .Y(_00178_));
 sky130_fd_sc_hd__nand2_1 _16656_ (.A(net251),
    .B(_05756_),
    .Y(_05789_));
 sky130_fd_sc_hd__o21ai_0 _16657_ (.A1(_05020_),
    .A2(_05756_),
    .B1(_05789_),
    .Y(_00179_));
 sky130_fd_sc_hd__nand2_1 _16658_ (.A(net250),
    .B(_05756_),
    .Y(_05790_));
 sky130_fd_sc_hd__o21ai_0 _16659_ (.A1(_05029_),
    .A2(_05756_),
    .B1(_05790_),
    .Y(_00180_));
 sky130_fd_sc_hd__nand2_1 _16660_ (.A(net249),
    .B(_05756_),
    .Y(_05791_));
 sky130_fd_sc_hd__o21ai_0 _16661_ (.A1(_05035_),
    .A2(_05756_),
    .B1(_05791_),
    .Y(_00181_));
 sky130_fd_sc_hd__nand2_1 _16662_ (.A(net248),
    .B(_05756_),
    .Y(_05792_));
 sky130_fd_sc_hd__o21ai_0 _16663_ (.A1(_05044_),
    .A2(_05756_),
    .B1(_05792_),
    .Y(_00182_));
 sky130_fd_sc_hd__nand2_1 _16664_ (.A(net247),
    .B(_05756_),
    .Y(_05793_));
 sky130_fd_sc_hd__o21ai_0 _16665_ (.A1(_05060_),
    .A2(_05756_),
    .B1(_05793_),
    .Y(_00184_));
 sky130_fd_sc_hd__mux2i_1 _16666_ (.A0(_05113_),
    .A1(net246),
    .S(_05756_),
    .Y(_05794_));
 sky130_fd_sc_hd__o21ai_0 _16667_ (.A1(_05112_),
    .A2(_05756_),
    .B1(_05794_),
    .Y(_00185_));
 sky130_fd_sc_hd__nand2_8 _16668_ (.A(_09784_),
    .B(_05474_),
    .Y(_05795_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1243 ();
 sky130_fd_sc_hd__nand2_1 _16671_ (.A(net582),
    .B(_05795_),
    .Y(_05798_));
 sky130_fd_sc_hd__o21ai_0 _16672_ (.A1(_05118_),
    .A2(_05795_),
    .B1(_05798_),
    .Y(_00193_));
 sky130_fd_sc_hd__nand2_1 _16673_ (.A(net581),
    .B(_05795_),
    .Y(_05799_));
 sky130_fd_sc_hd__o21ai_0 _16674_ (.A1(_05122_),
    .A2(_05795_),
    .B1(_05799_),
    .Y(_00204_));
 sky130_fd_sc_hd__nand2_1 _16675_ (.A(net580),
    .B(_05795_),
    .Y(_05800_));
 sky130_fd_sc_hd__o21ai_0 _16676_ (.A1(_05126_),
    .A2(_05795_),
    .B1(_05800_),
    .Y(_00215_));
 sky130_fd_sc_hd__nand2_1 _16677_ (.A(net579),
    .B(_05795_),
    .Y(_05801_));
 sky130_fd_sc_hd__o21ai_0 _16678_ (.A1(_05132_),
    .A2(_05795_),
    .B1(_05801_),
    .Y(_00218_));
 sky130_fd_sc_hd__nand2_1 _16679_ (.A(net577),
    .B(_05795_),
    .Y(_05802_));
 sky130_fd_sc_hd__o21ai_0 _16680_ (.A1(_05140_),
    .A2(_05795_),
    .B1(_05802_),
    .Y(_00219_));
 sky130_fd_sc_hd__nand2_1 _16681_ (.A(net576),
    .B(_05795_),
    .Y(_05803_));
 sky130_fd_sc_hd__o21ai_0 _16682_ (.A1(_05149_),
    .A2(_05795_),
    .B1(_05803_),
    .Y(_00220_));
 sky130_fd_sc_hd__nand2_1 _16683_ (.A(net575),
    .B(_05795_),
    .Y(_05804_));
 sky130_fd_sc_hd__o21ai_0 _16684_ (.A1(_05157_),
    .A2(_05795_),
    .B1(_05804_),
    .Y(_00221_));
 sky130_fd_sc_hd__nand2_1 _16685_ (.A(net574),
    .B(_05795_),
    .Y(_05805_));
 sky130_fd_sc_hd__o21ai_0 _16686_ (.A1(_05166_),
    .A2(_05795_),
    .B1(_05805_),
    .Y(_00222_));
 sky130_fd_sc_hd__nand2_1 _16687_ (.A(net573),
    .B(_05795_),
    .Y(_05806_));
 sky130_fd_sc_hd__o21ai_0 _16688_ (.A1(_05173_),
    .A2(_05795_),
    .B1(_05806_),
    .Y(_00223_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1242 ();
 sky130_fd_sc_hd__nand2_2 _16690_ (.A(net572),
    .B(_05795_),
    .Y(_05808_));
 sky130_fd_sc_hd__o21ai_0 _16691_ (.A1(_05183_),
    .A2(_05795_),
    .B1(_05808_),
    .Y(_00224_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1241 ();
 sky130_fd_sc_hd__nand2_1 _16693_ (.A(net571),
    .B(_05795_),
    .Y(_05810_));
 sky130_fd_sc_hd__o21ai_0 _16694_ (.A1(_05192_),
    .A2(_05795_),
    .B1(_05810_),
    .Y(_00194_));
 sky130_fd_sc_hd__nand2_1 _16695_ (.A(net570),
    .B(_05795_),
    .Y(_05811_));
 sky130_fd_sc_hd__o21ai_0 _16696_ (.A1(_05204_),
    .A2(_05795_),
    .B1(_05811_),
    .Y(_00195_));
 sky130_fd_sc_hd__nand2_1 _16697_ (.A(net569),
    .B(_05795_),
    .Y(_05812_));
 sky130_fd_sc_hd__o21ai_0 _16698_ (.A1(_05214_),
    .A2(_05795_),
    .B1(_05812_),
    .Y(_00196_));
 sky130_fd_sc_hd__nand2_1 _16699_ (.A(net568),
    .B(_05795_),
    .Y(_05813_));
 sky130_fd_sc_hd__o21ai_0 _16700_ (.A1(_05221_),
    .A2(_05795_),
    .B1(_05813_),
    .Y(_00197_));
 sky130_fd_sc_hd__nand2_1 _16701_ (.A(net566),
    .B(_05795_),
    .Y(_05814_));
 sky130_fd_sc_hd__o21ai_0 _16702_ (.A1(_05228_),
    .A2(_05795_),
    .B1(_05814_),
    .Y(_00198_));
 sky130_fd_sc_hd__nand2_1 _16703_ (.A(net565),
    .B(_05795_),
    .Y(_05815_));
 sky130_fd_sc_hd__o21ai_0 _16704_ (.A1(_05238_),
    .A2(_05795_),
    .B1(_05815_),
    .Y(_00199_));
 sky130_fd_sc_hd__nand2_1 _16705_ (.A(net564),
    .B(_05795_),
    .Y(_05816_));
 sky130_fd_sc_hd__o21ai_0 _16706_ (.A1(_05247_),
    .A2(_05795_),
    .B1(_05816_),
    .Y(_00200_));
 sky130_fd_sc_hd__nand2_1 _16707_ (.A(net563),
    .B(_05795_),
    .Y(_05817_));
 sky130_fd_sc_hd__o21ai_0 _16708_ (.A1(_05258_),
    .A2(_05795_),
    .B1(_05817_),
    .Y(_00201_));
 sky130_fd_sc_hd__nand2_1 _16709_ (.A(net562),
    .B(_05795_),
    .Y(_05818_));
 sky130_fd_sc_hd__o21ai_0 _16710_ (.A1(_05267_),
    .A2(_05795_),
    .B1(_05818_),
    .Y(_00202_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1240 ();
 sky130_fd_sc_hd__nand2_1 _16712_ (.A(net561),
    .B(_05795_),
    .Y(_05820_));
 sky130_fd_sc_hd__o21ai_0 _16713_ (.A1(_05280_),
    .A2(_05795_),
    .B1(_05820_),
    .Y(_00203_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1239 ();
 sky130_fd_sc_hd__nand2_1 _16715_ (.A(net560),
    .B(_05795_),
    .Y(_05822_));
 sky130_fd_sc_hd__o21ai_0 _16716_ (.A1(_05291_),
    .A2(_05795_),
    .B1(_05822_),
    .Y(_00205_));
 sky130_fd_sc_hd__nand2_1 _16717_ (.A(net559),
    .B(_05795_),
    .Y(_05823_));
 sky130_fd_sc_hd__o21ai_0 _16718_ (.A1(_05301_),
    .A2(_05795_),
    .B1(_05823_),
    .Y(_00206_));
 sky130_fd_sc_hd__nand2_1 _16719_ (.A(net558),
    .B(_05795_),
    .Y(_05824_));
 sky130_fd_sc_hd__o21ai_0 _16720_ (.A1(_05309_),
    .A2(_05795_),
    .B1(_05824_),
    .Y(_00207_));
 sky130_fd_sc_hd__nand2_1 _16721_ (.A(net557),
    .B(_05795_),
    .Y(_05825_));
 sky130_fd_sc_hd__o21ai_0 _16722_ (.A1(_05320_),
    .A2(_05795_),
    .B1(_05825_),
    .Y(_00208_));
 sky130_fd_sc_hd__nand2_1 _16723_ (.A(net555),
    .B(_05795_),
    .Y(_05826_));
 sky130_fd_sc_hd__o21ai_0 _16724_ (.A1(net1145),
    .A2(_05795_),
    .B1(_05826_),
    .Y(_00209_));
 sky130_fd_sc_hd__nand2_1 _16725_ (.A(net554),
    .B(_05795_),
    .Y(_05827_));
 sky130_fd_sc_hd__o21ai_0 _16726_ (.A1(_05339_),
    .A2(_05795_),
    .B1(_05827_),
    .Y(_00210_));
 sky130_fd_sc_hd__nand2_1 _16727_ (.A(net553),
    .B(_05795_),
    .Y(_05828_));
 sky130_fd_sc_hd__o21ai_0 _16728_ (.A1(_05347_),
    .A2(_05795_),
    .B1(_05828_),
    .Y(_00211_));
 sky130_fd_sc_hd__nand2_1 _16729_ (.A(net552),
    .B(_05795_),
    .Y(_05829_));
 sky130_fd_sc_hd__o21ai_0 _16730_ (.A1(_05358_),
    .A2(_05795_),
    .B1(_05829_),
    .Y(_00212_));
 sky130_fd_sc_hd__nand2_1 _16731_ (.A(net284),
    .B(_05795_),
    .Y(_05830_));
 sky130_fd_sc_hd__o21ai_0 _16732_ (.A1(_05372_),
    .A2(_05795_),
    .B1(_05830_),
    .Y(_00213_));
 sky130_fd_sc_hd__nand2_1 _16733_ (.A(net283),
    .B(_05795_),
    .Y(_05831_));
 sky130_fd_sc_hd__o21ai_0 _16734_ (.A1(_05380_),
    .A2(_05795_),
    .B1(_05831_),
    .Y(_00214_));
 sky130_fd_sc_hd__a21oi_1 _16735_ (.A1(_09784_),
    .A2(_05474_),
    .B1(net282),
    .Y(_05832_));
 sky130_fd_sc_hd__a31oi_1 _16736_ (.A1(_09784_),
    .A2(net1143),
    .A3(_05474_),
    .B1(_05832_),
    .Y(_00216_));
 sky130_fd_sc_hd__nand2_1 _16737_ (.A(net281),
    .B(_05795_),
    .Y(_05833_));
 sky130_fd_sc_hd__o21ai_0 _16738_ (.A1(_05430_),
    .A2(_05795_),
    .B1(_05833_),
    .Y(_00217_));
 sky130_fd_sc_hd__nand2_8 _16739_ (.A(_09739_),
    .B(_05516_),
    .Y(_05834_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1237 ();
 sky130_fd_sc_hd__nand2_1 _16742_ (.A(net618),
    .B(_05834_),
    .Y(_05837_));
 sky130_fd_sc_hd__o21ai_0 _16743_ (.A1(_04790_),
    .A2(_05834_),
    .B1(_05837_),
    .Y(_00225_));
 sky130_fd_sc_hd__nand2_1 _16744_ (.A(net617),
    .B(_05834_),
    .Y(_05838_));
 sky130_fd_sc_hd__o21ai_0 _16745_ (.A1(_04794_),
    .A2(_05834_),
    .B1(_05838_),
    .Y(_00236_));
 sky130_fd_sc_hd__nand2_1 _16746_ (.A(net616),
    .B(_05834_),
    .Y(_05839_));
 sky130_fd_sc_hd__o21ai_0 _16747_ (.A1(_04801_),
    .A2(_05834_),
    .B1(_05839_),
    .Y(_00247_));
 sky130_fd_sc_hd__nand2_1 _16748_ (.A(net615),
    .B(_05834_),
    .Y(_05840_));
 sky130_fd_sc_hd__o21ai_0 _16749_ (.A1(_04808_),
    .A2(_05834_),
    .B1(_05840_),
    .Y(_00250_));
 sky130_fd_sc_hd__nand2_1 _16750_ (.A(net614),
    .B(_05834_),
    .Y(_05841_));
 sky130_fd_sc_hd__o21ai_0 _16751_ (.A1(_04817_),
    .A2(_05834_),
    .B1(_05841_),
    .Y(_00251_));
 sky130_fd_sc_hd__nand2_1 _16752_ (.A(net613),
    .B(_05834_),
    .Y(_05842_));
 sky130_fd_sc_hd__o21ai_0 _16753_ (.A1(_04826_),
    .A2(_05834_),
    .B1(_05842_),
    .Y(_00252_));
 sky130_fd_sc_hd__nand2_1 _16754_ (.A(net611),
    .B(_05834_),
    .Y(_05843_));
 sky130_fd_sc_hd__o21ai_0 _16755_ (.A1(_04834_),
    .A2(_05834_),
    .B1(_05843_),
    .Y(_00253_));
 sky130_fd_sc_hd__nand2_1 _16756_ (.A(net610),
    .B(_05834_),
    .Y(_05844_));
 sky130_fd_sc_hd__o21ai_0 _16757_ (.A1(_04843_),
    .A2(_05834_),
    .B1(_05844_),
    .Y(_00254_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1236 ();
 sky130_fd_sc_hd__nand2_1 _16759_ (.A(net609),
    .B(_05834_),
    .Y(_05846_));
 sky130_fd_sc_hd__o21ai_0 _16760_ (.A1(_04852_),
    .A2(_05834_),
    .B1(_05846_),
    .Y(_00255_));
 sky130_fd_sc_hd__nand2_1 _16761_ (.A(net608),
    .B(_05834_),
    .Y(_05847_));
 sky130_fd_sc_hd__o21ai_0 _16762_ (.A1(_04860_),
    .A2(_05834_),
    .B1(_05847_),
    .Y(_00256_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1235 ();
 sky130_fd_sc_hd__nand2_1 _16764_ (.A(net607),
    .B(_05834_),
    .Y(_05849_));
 sky130_fd_sc_hd__o21ai_0 _16765_ (.A1(_04871_),
    .A2(_05834_),
    .B1(_05849_),
    .Y(_00226_));
 sky130_fd_sc_hd__nand2_1 _16766_ (.A(net606),
    .B(_05834_),
    .Y(_05850_));
 sky130_fd_sc_hd__o21ai_0 _16767_ (.A1(_04883_),
    .A2(_05834_),
    .B1(_05850_),
    .Y(_00227_));
 sky130_fd_sc_hd__nand2_1 _16768_ (.A(net605),
    .B(_05834_),
    .Y(_05851_));
 sky130_fd_sc_hd__o21ai_0 _16769_ (.A1(_04892_),
    .A2(_05834_),
    .B1(_05851_),
    .Y(_00228_));
 sky130_fd_sc_hd__nand2_1 _16770_ (.A(net604),
    .B(_05834_),
    .Y(_05852_));
 sky130_fd_sc_hd__o21ai_0 _16771_ (.A1(_04899_),
    .A2(_05834_),
    .B1(_05852_),
    .Y(_00229_));
 sky130_fd_sc_hd__nand2_1 _16772_ (.A(net603),
    .B(_05834_),
    .Y(_05853_));
 sky130_fd_sc_hd__o21ai_0 _16773_ (.A1(_04906_),
    .A2(_05834_),
    .B1(_05853_),
    .Y(_00230_));
 sky130_fd_sc_hd__nand2_1 _16774_ (.A(net602),
    .B(_05834_),
    .Y(_05854_));
 sky130_fd_sc_hd__o21ai_0 _16775_ (.A1(_04913_),
    .A2(_05834_),
    .B1(_05854_),
    .Y(_00231_));
 sky130_fd_sc_hd__nand2_1 _16776_ (.A(net599),
    .B(_05834_),
    .Y(_05855_));
 sky130_fd_sc_hd__o21ai_0 _16777_ (.A1(_04923_),
    .A2(_05834_),
    .B1(_05855_),
    .Y(_00232_));
 sky130_fd_sc_hd__nand2_1 _16778_ (.A(net598),
    .B(_05834_),
    .Y(_05856_));
 sky130_fd_sc_hd__o21ai_0 _16779_ (.A1(_04932_),
    .A2(_05834_),
    .B1(_05856_),
    .Y(_00233_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1234 ();
 sky130_fd_sc_hd__nand2_1 _16781_ (.A(net597),
    .B(_05834_),
    .Y(_05858_));
 sky130_fd_sc_hd__o21ai_0 _16782_ (.A1(_04939_),
    .A2(_05834_),
    .B1(_05858_),
    .Y(_00234_));
 sky130_fd_sc_hd__nand2_1 _16783_ (.A(net596),
    .B(_05834_),
    .Y(_05859_));
 sky130_fd_sc_hd__o21ai_0 _16784_ (.A1(_04951_),
    .A2(_05834_),
    .B1(_05859_),
    .Y(_00235_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1233 ();
 sky130_fd_sc_hd__nand2_1 _16786_ (.A(net595),
    .B(_05834_),
    .Y(_05861_));
 sky130_fd_sc_hd__o21ai_0 _16787_ (.A1(_04960_),
    .A2(_05834_),
    .B1(_05861_),
    .Y(_00237_));
 sky130_fd_sc_hd__nand2_1 _16788_ (.A(net594),
    .B(_05834_),
    .Y(_05862_));
 sky130_fd_sc_hd__o21ai_0 _16789_ (.A1(_04974_),
    .A2(_05834_),
    .B1(_05862_),
    .Y(_00238_));
 sky130_fd_sc_hd__nand2_1 _16790_ (.A(net593),
    .B(_05834_),
    .Y(_05863_));
 sky130_fd_sc_hd__o21ai_0 _16791_ (.A1(_04984_),
    .A2(_05834_),
    .B1(_05863_),
    .Y(_00239_));
 sky130_fd_sc_hd__nand2_1 _16792_ (.A(net592),
    .B(_05834_),
    .Y(_05864_));
 sky130_fd_sc_hd__o21ai_0 _16793_ (.A1(_04990_),
    .A2(_05834_),
    .B1(_05864_),
    .Y(_00240_));
 sky130_fd_sc_hd__nand2_1 _16794_ (.A(net591),
    .B(_05834_),
    .Y(_05865_));
 sky130_fd_sc_hd__o21ai_0 _16795_ (.A1(net1129),
    .A2(_05834_),
    .B1(_05865_),
    .Y(_00241_));
 sky130_fd_sc_hd__nand2_1 _16796_ (.A(net590),
    .B(_05834_),
    .Y(_05866_));
 sky130_fd_sc_hd__o21ai_0 _16797_ (.A1(_05011_),
    .A2(_05834_),
    .B1(_05866_),
    .Y(_00242_));
 sky130_fd_sc_hd__nand2_1 _16798_ (.A(net588),
    .B(_05834_),
    .Y(_05867_));
 sky130_fd_sc_hd__o21ai_0 _16799_ (.A1(_05020_),
    .A2(_05834_),
    .B1(_05867_),
    .Y(_00243_));
 sky130_fd_sc_hd__nand2_1 _16800_ (.A(net587),
    .B(_05834_),
    .Y(_05868_));
 sky130_fd_sc_hd__o21ai_0 _16801_ (.A1(_05029_),
    .A2(_05834_),
    .B1(_05868_),
    .Y(_00244_));
 sky130_fd_sc_hd__nand2_1 _16802_ (.A(net586),
    .B(_05834_),
    .Y(_05869_));
 sky130_fd_sc_hd__o21ai_0 _16803_ (.A1(_05035_),
    .A2(_05834_),
    .B1(_05869_),
    .Y(_00245_));
 sky130_fd_sc_hd__nand2_1 _16804_ (.A(net585),
    .B(_05834_),
    .Y(_05870_));
 sky130_fd_sc_hd__o21ai_0 _16805_ (.A1(_05044_),
    .A2(_05834_),
    .B1(_05870_),
    .Y(_00246_));
 sky130_fd_sc_hd__nand2_1 _16806_ (.A(net584),
    .B(_05834_),
    .Y(_05871_));
 sky130_fd_sc_hd__o21ai_0 _16807_ (.A1(_05060_),
    .A2(_05834_),
    .B1(_05871_),
    .Y(_00248_));
 sky130_fd_sc_hd__mux2i_1 _16808_ (.A0(_05113_),
    .A1(net583),
    .S(_05834_),
    .Y(_05872_));
 sky130_fd_sc_hd__o21ai_0 _16809_ (.A1(_05112_),
    .A2(_05834_),
    .B1(_05872_),
    .Y(_00249_));
 sky130_fd_sc_hd__nand2_8 _16810_ (.A(net551),
    .B(_05557_),
    .Y(_05873_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1231 ();
 sky130_fd_sc_hd__nand2_1 _16813_ (.A(net653),
    .B(_05873_),
    .Y(_05876_));
 sky130_fd_sc_hd__o21ai_0 _16814_ (.A1(_05118_),
    .A2(_05873_),
    .B1(_05876_),
    .Y(_00257_));
 sky130_fd_sc_hd__nand2_1 _16815_ (.A(net652),
    .B(_05873_),
    .Y(_05877_));
 sky130_fd_sc_hd__o21ai_0 _16816_ (.A1(_05122_),
    .A2(_05873_),
    .B1(_05877_),
    .Y(_00268_));
 sky130_fd_sc_hd__nand2_1 _16817_ (.A(net651),
    .B(_05873_),
    .Y(_05878_));
 sky130_fd_sc_hd__o21ai_0 _16818_ (.A1(_05126_),
    .A2(_05873_),
    .B1(_05878_),
    .Y(_00279_));
 sky130_fd_sc_hd__nand2_1 _16819_ (.A(net650),
    .B(_05873_),
    .Y(_05879_));
 sky130_fd_sc_hd__o21ai_0 _16820_ (.A1(_05132_),
    .A2(_05873_),
    .B1(_05879_),
    .Y(_00282_));
 sky130_fd_sc_hd__nand2_1 _16821_ (.A(net649),
    .B(_05873_),
    .Y(_05880_));
 sky130_fd_sc_hd__o21ai_0 _16822_ (.A1(_05140_),
    .A2(_05873_),
    .B1(_05880_),
    .Y(_00283_));
 sky130_fd_sc_hd__nand2_1 _16823_ (.A(net648),
    .B(_05873_),
    .Y(_05881_));
 sky130_fd_sc_hd__o21ai_0 _16824_ (.A1(_05149_),
    .A2(_05873_),
    .B1(_05881_),
    .Y(_00284_));
 sky130_fd_sc_hd__nand2_1 _16825_ (.A(net647),
    .B(_05873_),
    .Y(_05882_));
 sky130_fd_sc_hd__o21ai_0 _16826_ (.A1(_05157_),
    .A2(_05873_),
    .B1(_05882_),
    .Y(_00285_));
 sky130_fd_sc_hd__nand2_1 _16827_ (.A(net646),
    .B(_05873_),
    .Y(_05883_));
 sky130_fd_sc_hd__o21ai_0 _16828_ (.A1(_05166_),
    .A2(_05873_),
    .B1(_05883_),
    .Y(_00286_));
 sky130_fd_sc_hd__nand2_1 _16829_ (.A(net644),
    .B(_05873_),
    .Y(_05884_));
 sky130_fd_sc_hd__o21ai_0 _16830_ (.A1(_05173_),
    .A2(_05873_),
    .B1(_05884_),
    .Y(_00287_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1230 ();
 sky130_fd_sc_hd__nand2_1 _16832_ (.A(net643),
    .B(_05873_),
    .Y(_05886_));
 sky130_fd_sc_hd__o21ai_0 _16833_ (.A1(_05183_),
    .A2(_05873_),
    .B1(_05886_),
    .Y(_00288_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1229 ();
 sky130_fd_sc_hd__nand2_1 _16835_ (.A(net642),
    .B(_05873_),
    .Y(_05888_));
 sky130_fd_sc_hd__o21ai_0 _16836_ (.A1(_05192_),
    .A2(_05873_),
    .B1(_05888_),
    .Y(_00258_));
 sky130_fd_sc_hd__nand2_1 _16837_ (.A(net641),
    .B(_05873_),
    .Y(_05889_));
 sky130_fd_sc_hd__o21ai_0 _16838_ (.A1(_05204_),
    .A2(_05873_),
    .B1(_05889_),
    .Y(_00259_));
 sky130_fd_sc_hd__nand2_1 _16839_ (.A(net640),
    .B(_05873_),
    .Y(_05890_));
 sky130_fd_sc_hd__o21ai_0 _16840_ (.A1(_05214_),
    .A2(_05873_),
    .B1(_05890_),
    .Y(_00260_));
 sky130_fd_sc_hd__nand2_1 _16841_ (.A(net639),
    .B(_05873_),
    .Y(_05891_));
 sky130_fd_sc_hd__o21ai_0 _16842_ (.A1(_05221_),
    .A2(_05873_),
    .B1(_05891_),
    .Y(_00261_));
 sky130_fd_sc_hd__nand2_1 _16843_ (.A(net638),
    .B(_05873_),
    .Y(_05892_));
 sky130_fd_sc_hd__o21ai_0 _16844_ (.A1(_05228_),
    .A2(_05873_),
    .B1(_05892_),
    .Y(_00262_));
 sky130_fd_sc_hd__nand2_1 _16845_ (.A(net637),
    .B(_05873_),
    .Y(_05893_));
 sky130_fd_sc_hd__o21ai_0 _16846_ (.A1(_05238_),
    .A2(_05873_),
    .B1(_05893_),
    .Y(_00263_));
 sky130_fd_sc_hd__nand2_1 _16847_ (.A(net636),
    .B(_05873_),
    .Y(_05894_));
 sky130_fd_sc_hd__o21ai_0 _16848_ (.A1(_05247_),
    .A2(_05873_),
    .B1(_05894_),
    .Y(_00264_));
 sky130_fd_sc_hd__nand2_1 _16849_ (.A(net635),
    .B(_05873_),
    .Y(_05895_));
 sky130_fd_sc_hd__o21ai_0 _16850_ (.A1(_05258_),
    .A2(_05873_),
    .B1(_05895_),
    .Y(_00265_));
 sky130_fd_sc_hd__nand2_1 _16851_ (.A(net633),
    .B(_05873_),
    .Y(_05896_));
 sky130_fd_sc_hd__o21ai_0 _16852_ (.A1(_05267_),
    .A2(_05873_),
    .B1(_05896_),
    .Y(_00266_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1228 ();
 sky130_fd_sc_hd__nand2_1 _16854_ (.A(net632),
    .B(_05873_),
    .Y(_05898_));
 sky130_fd_sc_hd__o21ai_0 _16855_ (.A1(_05280_),
    .A2(_05873_),
    .B1(_05898_),
    .Y(_00267_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1227 ();
 sky130_fd_sc_hd__nand2_1 _16857_ (.A(net631),
    .B(_05873_),
    .Y(_05900_));
 sky130_fd_sc_hd__o21ai_0 _16858_ (.A1(_05291_),
    .A2(_05873_),
    .B1(_05900_),
    .Y(_00269_));
 sky130_fd_sc_hd__nand2_1 _16859_ (.A(net630),
    .B(_05873_),
    .Y(_05901_));
 sky130_fd_sc_hd__o21ai_0 _16860_ (.A1(_05301_),
    .A2(_05873_),
    .B1(_05901_),
    .Y(_00270_));
 sky130_fd_sc_hd__nand2_1 _16861_ (.A(net629),
    .B(_05873_),
    .Y(_05902_));
 sky130_fd_sc_hd__o21ai_0 _16862_ (.A1(_05309_),
    .A2(_05873_),
    .B1(_05902_),
    .Y(_00271_));
 sky130_fd_sc_hd__nand2_1 _16863_ (.A(net628),
    .B(_05873_),
    .Y(_05903_));
 sky130_fd_sc_hd__o21ai_0 _16864_ (.A1(_05320_),
    .A2(_05873_),
    .B1(_05903_),
    .Y(_00272_));
 sky130_fd_sc_hd__nand2_1 _16865_ (.A(net627),
    .B(_05873_),
    .Y(_05904_));
 sky130_fd_sc_hd__o21ai_0 _16866_ (.A1(net1145),
    .A2(_05873_),
    .B1(_05904_),
    .Y(_00273_));
 sky130_fd_sc_hd__nand2_1 _16867_ (.A(net626),
    .B(_05873_),
    .Y(_05905_));
 sky130_fd_sc_hd__o21ai_0 _16868_ (.A1(_05339_),
    .A2(_05873_),
    .B1(_05905_),
    .Y(_00274_));
 sky130_fd_sc_hd__nand2_1 _16869_ (.A(net625),
    .B(_05873_),
    .Y(_05906_));
 sky130_fd_sc_hd__o21ai_0 _16870_ (.A1(_05347_),
    .A2(_05873_),
    .B1(_05906_),
    .Y(_00275_));
 sky130_fd_sc_hd__nand2_1 _16871_ (.A(net624),
    .B(_05873_),
    .Y(_05907_));
 sky130_fd_sc_hd__o21ai_0 _16872_ (.A1(_05358_),
    .A2(_05873_),
    .B1(_05907_),
    .Y(_00276_));
 sky130_fd_sc_hd__nand2_1 _16873_ (.A(net622),
    .B(_05873_),
    .Y(_05908_));
 sky130_fd_sc_hd__o21ai_0 _16874_ (.A1(_05372_),
    .A2(_05873_),
    .B1(_05908_),
    .Y(_00277_));
 sky130_fd_sc_hd__nand2_1 _16875_ (.A(net621),
    .B(_05873_),
    .Y(_05909_));
 sky130_fd_sc_hd__o21ai_0 _16876_ (.A1(_05380_),
    .A2(_05873_),
    .B1(_05909_),
    .Y(_00278_));
 sky130_fd_sc_hd__a21oi_1 _16877_ (.A1(_09784_),
    .A2(_05557_),
    .B1(net620),
    .Y(_05910_));
 sky130_fd_sc_hd__a31oi_1 _16878_ (.A1(_09784_),
    .A2(net1143),
    .A3(_05557_),
    .B1(_05910_),
    .Y(_00280_));
 sky130_fd_sc_hd__nand2_1 _16879_ (.A(net619),
    .B(_05873_),
    .Y(_05911_));
 sky130_fd_sc_hd__o21ai_0 _16880_ (.A1(_05430_),
    .A2(_05873_),
    .B1(_05911_),
    .Y(_00281_));
 sky130_fd_sc_hd__nand2_8 _16881_ (.A(_09739_),
    .B(_05598_),
    .Y(_05912_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1225 ();
 sky130_fd_sc_hd__nand2_1 _16884_ (.A(net688),
    .B(_05912_),
    .Y(_05915_));
 sky130_fd_sc_hd__o21ai_0 _16885_ (.A1(_04790_),
    .A2(_05912_),
    .B1(_05915_),
    .Y(_00289_));
 sky130_fd_sc_hd__nand2_1 _16886_ (.A(net687),
    .B(_05912_),
    .Y(_05916_));
 sky130_fd_sc_hd__o21ai_0 _16887_ (.A1(_04794_),
    .A2(_05912_),
    .B1(_05916_),
    .Y(_00300_));
 sky130_fd_sc_hd__nand2_1 _16888_ (.A(net686),
    .B(_05912_),
    .Y(_05917_));
 sky130_fd_sc_hd__o21ai_0 _16889_ (.A1(_04801_),
    .A2(_05912_),
    .B1(_05917_),
    .Y(_00311_));
 sky130_fd_sc_hd__nand2_1 _16890_ (.A(net685),
    .B(_05912_),
    .Y(_05918_));
 sky130_fd_sc_hd__o21ai_0 _16891_ (.A1(_04808_),
    .A2(_05912_),
    .B1(_05918_),
    .Y(_00314_));
 sky130_fd_sc_hd__nand2_1 _16892_ (.A(net684),
    .B(_05912_),
    .Y(_05919_));
 sky130_fd_sc_hd__o21ai_0 _16893_ (.A1(_04817_),
    .A2(_05912_),
    .B1(_05919_),
    .Y(_00315_));
 sky130_fd_sc_hd__nand2_1 _16894_ (.A(net683),
    .B(_05912_),
    .Y(_05920_));
 sky130_fd_sc_hd__o21ai_0 _16895_ (.A1(_04826_),
    .A2(_05912_),
    .B1(_05920_),
    .Y(_00316_));
 sky130_fd_sc_hd__nand2_1 _16896_ (.A(net682),
    .B(_05912_),
    .Y(_05921_));
 sky130_fd_sc_hd__o21ai_0 _16897_ (.A1(_04834_),
    .A2(_05912_),
    .B1(_05921_),
    .Y(_00317_));
 sky130_fd_sc_hd__nand2_1 _16898_ (.A(net681),
    .B(_05912_),
    .Y(_05922_));
 sky130_fd_sc_hd__o21ai_0 _16899_ (.A1(_04843_),
    .A2(_05912_),
    .B1(_05922_),
    .Y(_00318_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1224 ();
 sky130_fd_sc_hd__nand2_1 _16901_ (.A(net680),
    .B(_05912_),
    .Y(_05924_));
 sky130_fd_sc_hd__o21ai_0 _16902_ (.A1(_04852_),
    .A2(_05912_),
    .B1(_05924_),
    .Y(_00319_));
 sky130_fd_sc_hd__nand2_1 _16903_ (.A(net679),
    .B(_05912_),
    .Y(_05925_));
 sky130_fd_sc_hd__o21ai_0 _16904_ (.A1(_04860_),
    .A2(_05912_),
    .B1(_05925_),
    .Y(_00320_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1223 ();
 sky130_fd_sc_hd__nand2_1 _16906_ (.A(net677),
    .B(_05912_),
    .Y(_05927_));
 sky130_fd_sc_hd__o21ai_0 _16907_ (.A1(_04871_),
    .A2(_05912_),
    .B1(_05927_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_1 _16908_ (.A(net676),
    .B(_05912_),
    .Y(_05928_));
 sky130_fd_sc_hd__o21ai_0 _16909_ (.A1(_04883_),
    .A2(_05912_),
    .B1(_05928_),
    .Y(_00291_));
 sky130_fd_sc_hd__nand2_1 _16910_ (.A(net675),
    .B(_05912_),
    .Y(_05929_));
 sky130_fd_sc_hd__o21ai_0 _16911_ (.A1(_04892_),
    .A2(_05912_),
    .B1(_05929_),
    .Y(_00292_));
 sky130_fd_sc_hd__nand2_1 _16912_ (.A(net674),
    .B(_05912_),
    .Y(_05930_));
 sky130_fd_sc_hd__o21ai_0 _16913_ (.A1(_04899_),
    .A2(_05912_),
    .B1(_05930_),
    .Y(_00293_));
 sky130_fd_sc_hd__nand2_1 _16914_ (.A(net673),
    .B(_05912_),
    .Y(_05931_));
 sky130_fd_sc_hd__o21ai_0 _16915_ (.A1(_04906_),
    .A2(_05912_),
    .B1(_05931_),
    .Y(_00294_));
 sky130_fd_sc_hd__nand2_1 _16916_ (.A(net672),
    .B(_05912_),
    .Y(_05932_));
 sky130_fd_sc_hd__o21ai_0 _16917_ (.A1(_04913_),
    .A2(_05912_),
    .B1(_05932_),
    .Y(_00295_));
 sky130_fd_sc_hd__nand2_1 _16918_ (.A(net671),
    .B(_05912_),
    .Y(_05933_));
 sky130_fd_sc_hd__o21ai_0 _16919_ (.A1(_04923_),
    .A2(_05912_),
    .B1(_05933_),
    .Y(_00296_));
 sky130_fd_sc_hd__nand2_1 _16920_ (.A(net670),
    .B(_05912_),
    .Y(_05934_));
 sky130_fd_sc_hd__o21ai_0 _16921_ (.A1(_04932_),
    .A2(_05912_),
    .B1(_05934_),
    .Y(_00297_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1222 ();
 sky130_fd_sc_hd__nand2_1 _16923_ (.A(net669),
    .B(_05912_),
    .Y(_05936_));
 sky130_fd_sc_hd__o21ai_0 _16924_ (.A1(_04939_),
    .A2(_05912_),
    .B1(_05936_),
    .Y(_00298_));
 sky130_fd_sc_hd__nand2_1 _16925_ (.A(net668),
    .B(_05912_),
    .Y(_05937_));
 sky130_fd_sc_hd__o21ai_0 _16926_ (.A1(_04951_),
    .A2(_05912_),
    .B1(_05937_),
    .Y(_00299_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1221 ();
 sky130_fd_sc_hd__nand2_2 _16928_ (.A(net666),
    .B(_05912_),
    .Y(_05939_));
 sky130_fd_sc_hd__o21ai_0 _16929_ (.A1(_04960_),
    .A2(_05912_),
    .B1(_05939_),
    .Y(_00301_));
 sky130_fd_sc_hd__nand2_1 _16930_ (.A(net665),
    .B(_05912_),
    .Y(_05940_));
 sky130_fd_sc_hd__o21ai_0 _16931_ (.A1(_04974_),
    .A2(_05912_),
    .B1(_05940_),
    .Y(_00302_));
 sky130_fd_sc_hd__nand2_1 _16932_ (.A(net664),
    .B(_05912_),
    .Y(_05941_));
 sky130_fd_sc_hd__o21ai_0 _16933_ (.A1(_04984_),
    .A2(_05912_),
    .B1(_05941_),
    .Y(_00303_));
 sky130_fd_sc_hd__nand2_1 _16934_ (.A(net663),
    .B(_05912_),
    .Y(_05942_));
 sky130_fd_sc_hd__o21ai_0 _16935_ (.A1(_04990_),
    .A2(_05912_),
    .B1(_05942_),
    .Y(_00304_));
 sky130_fd_sc_hd__nand2_1 _16936_ (.A(net662),
    .B(_05912_),
    .Y(_05943_));
 sky130_fd_sc_hd__o21ai_0 _16937_ (.A1(net1129),
    .A2(_05912_),
    .B1(_05943_),
    .Y(_00305_));
 sky130_fd_sc_hd__nand2_1 _16938_ (.A(net661),
    .B(_05912_),
    .Y(_05944_));
 sky130_fd_sc_hd__o21ai_0 _16939_ (.A1(_05011_),
    .A2(_05912_),
    .B1(_05944_),
    .Y(_00306_));
 sky130_fd_sc_hd__nand2_1 _16940_ (.A(net660),
    .B(_05912_),
    .Y(_05945_));
 sky130_fd_sc_hd__o21ai_0 _16941_ (.A1(_05020_),
    .A2(_05912_),
    .B1(_05945_),
    .Y(_00307_));
 sky130_fd_sc_hd__nand2_1 _16942_ (.A(net659),
    .B(_05912_),
    .Y(_05946_));
 sky130_fd_sc_hd__o21ai_0 _16943_ (.A1(_05029_),
    .A2(_05912_),
    .B1(_05946_),
    .Y(_00308_));
 sky130_fd_sc_hd__nand2_1 _16944_ (.A(net658),
    .B(_05912_),
    .Y(_05947_));
 sky130_fd_sc_hd__o21ai_0 _16945_ (.A1(_05035_),
    .A2(_05912_),
    .B1(_05947_),
    .Y(_00309_));
 sky130_fd_sc_hd__nand2_1 _16946_ (.A(net657),
    .B(_05912_),
    .Y(_05948_));
 sky130_fd_sc_hd__o21ai_0 _16947_ (.A1(_05044_),
    .A2(_05912_),
    .B1(_05948_),
    .Y(_00310_));
 sky130_fd_sc_hd__nand2_1 _16948_ (.A(net655),
    .B(_05912_),
    .Y(_05949_));
 sky130_fd_sc_hd__o21ai_0 _16949_ (.A1(_05060_),
    .A2(_05912_),
    .B1(_05949_),
    .Y(_00312_));
 sky130_fd_sc_hd__mux2i_1 _16950_ (.A0(_05113_),
    .A1(net654),
    .S(_05912_),
    .Y(_05950_));
 sky130_fd_sc_hd__o21ai_0 _16951_ (.A1(_05112_),
    .A2(_05912_),
    .B1(_05950_),
    .Y(_00313_));
 sky130_fd_sc_hd__nor2b_4 _16952_ (.A(net1039),
    .B_N(_13541_),
    .Y(_05951_));
 sky130_fd_sc_hd__nand2_8 _16953_ (.A(net551),
    .B(_05951_),
    .Y(_05952_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1219 ();
 sky130_fd_sc_hd__nand2_1 _16956_ (.A(net725),
    .B(_05952_),
    .Y(_05955_));
 sky130_fd_sc_hd__o21ai_0 _16957_ (.A1(_05118_),
    .A2(_05952_),
    .B1(_05955_),
    .Y(_00321_));
 sky130_fd_sc_hd__nand2_1 _16958_ (.A(net724),
    .B(_05952_),
    .Y(_05956_));
 sky130_fd_sc_hd__o21ai_0 _16959_ (.A1(_05122_),
    .A2(_05952_),
    .B1(_05956_),
    .Y(_00332_));
 sky130_fd_sc_hd__nand2_1 _16960_ (.A(net722),
    .B(_05952_),
    .Y(_05957_));
 sky130_fd_sc_hd__o21ai_0 _16961_ (.A1(_05126_),
    .A2(_05952_),
    .B1(_05957_),
    .Y(_00343_));
 sky130_fd_sc_hd__nand2_1 _16962_ (.A(net721),
    .B(_05952_),
    .Y(_05958_));
 sky130_fd_sc_hd__o21ai_0 _16963_ (.A1(_05132_),
    .A2(_05952_),
    .B1(_05958_),
    .Y(_00346_));
 sky130_fd_sc_hd__nand2_1 _16964_ (.A(net720),
    .B(_05952_),
    .Y(_05959_));
 sky130_fd_sc_hd__o21ai_0 _16965_ (.A1(_05140_),
    .A2(_05952_),
    .B1(_05959_),
    .Y(_00347_));
 sky130_fd_sc_hd__nand2_1 _16966_ (.A(net719),
    .B(_05952_),
    .Y(_05960_));
 sky130_fd_sc_hd__o21ai_0 _16967_ (.A1(_05149_),
    .A2(_05952_),
    .B1(_05960_),
    .Y(_00348_));
 sky130_fd_sc_hd__nand2_1 _16968_ (.A(net718),
    .B(_05952_),
    .Y(_05961_));
 sky130_fd_sc_hd__o21ai_0 _16969_ (.A1(_05157_),
    .A2(_05952_),
    .B1(_05961_),
    .Y(_00349_));
 sky130_fd_sc_hd__nand2_1 _16970_ (.A(net717),
    .B(_05952_),
    .Y(_05962_));
 sky130_fd_sc_hd__o21ai_0 _16971_ (.A1(_05166_),
    .A2(_05952_),
    .B1(_05962_),
    .Y(_00350_));
 sky130_fd_sc_hd__nand2_1 _16972_ (.A(net716),
    .B(_05952_),
    .Y(_05963_));
 sky130_fd_sc_hd__o21ai_0 _16973_ (.A1(_05173_),
    .A2(_05952_),
    .B1(_05963_),
    .Y(_00351_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1218 ();
 sky130_fd_sc_hd__nand2_1 _16975_ (.A(net715),
    .B(_05952_),
    .Y(_05965_));
 sky130_fd_sc_hd__o21ai_0 _16976_ (.A1(_05183_),
    .A2(_05952_),
    .B1(_05965_),
    .Y(_00352_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1217 ();
 sky130_fd_sc_hd__nand2_1 _16978_ (.A(net714),
    .B(_05952_),
    .Y(_05967_));
 sky130_fd_sc_hd__o21ai_0 _16979_ (.A1(_05192_),
    .A2(_05952_),
    .B1(_05967_),
    .Y(_00322_));
 sky130_fd_sc_hd__nand2_1 _16980_ (.A(net713),
    .B(_05952_),
    .Y(_05968_));
 sky130_fd_sc_hd__o21ai_0 _16981_ (.A1(_05204_),
    .A2(_05952_),
    .B1(_05968_),
    .Y(_00323_));
 sky130_fd_sc_hd__nand2_1 _16982_ (.A(net710),
    .B(_05952_),
    .Y(_05969_));
 sky130_fd_sc_hd__o21ai_0 _16983_ (.A1(_05214_),
    .A2(_05952_),
    .B1(_05969_),
    .Y(_00324_));
 sky130_fd_sc_hd__nand2_1 _16984_ (.A(net709),
    .B(_05952_),
    .Y(_05970_));
 sky130_fd_sc_hd__o21ai_0 _16985_ (.A1(_05221_),
    .A2(_05952_),
    .B1(_05970_),
    .Y(_00325_));
 sky130_fd_sc_hd__nand2_1 _16986_ (.A(net708),
    .B(_05952_),
    .Y(_05971_));
 sky130_fd_sc_hd__o21ai_0 _16987_ (.A1(_05228_),
    .A2(_05952_),
    .B1(_05971_),
    .Y(_00326_));
 sky130_fd_sc_hd__nand2_1 _16988_ (.A(net707),
    .B(_05952_),
    .Y(_05972_));
 sky130_fd_sc_hd__o21ai_0 _16989_ (.A1(_05238_),
    .A2(_05952_),
    .B1(_05972_),
    .Y(_00327_));
 sky130_fd_sc_hd__nand2_1 _16990_ (.A(net706),
    .B(_05952_),
    .Y(_05973_));
 sky130_fd_sc_hd__o21ai_0 _16991_ (.A1(_05247_),
    .A2(_05952_),
    .B1(_05973_),
    .Y(_00328_));
 sky130_fd_sc_hd__nand2_1 _16992_ (.A(net705),
    .B(_05952_),
    .Y(_05974_));
 sky130_fd_sc_hd__o21ai_0 _16993_ (.A1(_05258_),
    .A2(_05952_),
    .B1(_05974_),
    .Y(_00329_));
 sky130_fd_sc_hd__nand2_1 _16994_ (.A(net704),
    .B(_05952_),
    .Y(_05975_));
 sky130_fd_sc_hd__o21ai_0 _16995_ (.A1(_05267_),
    .A2(_05952_),
    .B1(_05975_),
    .Y(_00330_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1216 ();
 sky130_fd_sc_hd__nand2_1 _16997_ (.A(net703),
    .B(_05952_),
    .Y(_05977_));
 sky130_fd_sc_hd__o21ai_0 _16998_ (.A1(_05280_),
    .A2(_05952_),
    .B1(_05977_),
    .Y(_00331_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1215 ();
 sky130_fd_sc_hd__nand2_1 _17000_ (.A(net702),
    .B(_05952_),
    .Y(_05979_));
 sky130_fd_sc_hd__o21ai_0 _17001_ (.A1(_05291_),
    .A2(_05952_),
    .B1(_05979_),
    .Y(_00333_));
 sky130_fd_sc_hd__nand2_1 _17002_ (.A(net701),
    .B(_05952_),
    .Y(_05980_));
 sky130_fd_sc_hd__o21ai_0 _17003_ (.A1(_05301_),
    .A2(_05952_),
    .B1(_05980_),
    .Y(_00334_));
 sky130_fd_sc_hd__nand2_1 _17004_ (.A(net699),
    .B(_05952_),
    .Y(_05981_));
 sky130_fd_sc_hd__o21ai_0 _17005_ (.A1(_05309_),
    .A2(_05952_),
    .B1(_05981_),
    .Y(_00335_));
 sky130_fd_sc_hd__nand2_1 _17006_ (.A(net698),
    .B(_05952_),
    .Y(_05982_));
 sky130_fd_sc_hd__o21ai_0 _17007_ (.A1(_05320_),
    .A2(_05952_),
    .B1(_05982_),
    .Y(_00336_));
 sky130_fd_sc_hd__nand2_1 _17008_ (.A(net697),
    .B(_05952_),
    .Y(_05983_));
 sky130_fd_sc_hd__o21ai_0 _17009_ (.A1(net1145),
    .A2(_05952_),
    .B1(_05983_),
    .Y(_00337_));
 sky130_fd_sc_hd__nand2_1 _17010_ (.A(net696),
    .B(_05952_),
    .Y(_05984_));
 sky130_fd_sc_hd__o21ai_0 _17011_ (.A1(_05339_),
    .A2(_05952_),
    .B1(_05984_),
    .Y(_00338_));
 sky130_fd_sc_hd__nand2_1 _17012_ (.A(net695),
    .B(_05952_),
    .Y(_05985_));
 sky130_fd_sc_hd__o21ai_0 _17013_ (.A1(_05347_),
    .A2(_05952_),
    .B1(_05985_),
    .Y(_00339_));
 sky130_fd_sc_hd__nand2_1 _17014_ (.A(net694),
    .B(_05952_),
    .Y(_05986_));
 sky130_fd_sc_hd__o21ai_0 _17015_ (.A1(_05358_),
    .A2(_05952_),
    .B1(_05986_),
    .Y(_00340_));
 sky130_fd_sc_hd__nand2_1 _17016_ (.A(net693),
    .B(_05952_),
    .Y(_05987_));
 sky130_fd_sc_hd__o21ai_0 _17017_ (.A1(_05372_),
    .A2(_05952_),
    .B1(_05987_),
    .Y(_00341_));
 sky130_fd_sc_hd__nand2_1 _17018_ (.A(net692),
    .B(_05952_),
    .Y(_05988_));
 sky130_fd_sc_hd__o21ai_0 _17019_ (.A1(_05380_),
    .A2(_05952_),
    .B1(_05988_),
    .Y(_00342_));
 sky130_fd_sc_hd__a21oi_1 _17020_ (.A1(net551),
    .A2(_05951_),
    .B1(net691),
    .Y(_05989_));
 sky130_fd_sc_hd__a31oi_1 _17021_ (.A1(net551),
    .A2(net1143),
    .A3(_05951_),
    .B1(_05989_),
    .Y(_00344_));
 sky130_fd_sc_hd__nand2_1 _17022_ (.A(net690),
    .B(_05952_),
    .Y(_05990_));
 sky130_fd_sc_hd__o21ai_0 _17023_ (.A1(_05430_),
    .A2(_05952_),
    .B1(_05990_),
    .Y(_00345_));
 sky130_fd_sc_hd__or2_4 _17024_ (.A(net343),
    .B(\hash.CA2.f_dash[0] ),
    .X(_12653_));
 sky130_fd_sc_hd__inv_1 _17025_ (.A(_12653_),
    .Y(_00875_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1214 ();
 sky130_fd_sc_hd__nor2_4 _17027_ (.A(net344),
    .B(\hash.CA2.e_dash[0] ),
    .Y(_00843_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1208 ();
 sky130_fd_sc_hd__clkinvlp_4 _17034_ (.A(_12109_),
    .Y(_05998_));
 sky130_fd_sc_hd__nor2_2 _17035_ (.A(net340),
    .B(_05998_),
    .Y(_05999_));
 sky130_fd_sc_hd__inv_1 _17036_ (.A(_05999_),
    .Y(\hash.CA1.S0.X[2] ));
 sky130_fd_sc_hd__xnor2_1 _17037_ (.A(_13544_),
    .B(_05999_),
    .Y(_00680_));
 sky130_fd_sc_hd__xor2_1 _17038_ (.A(_12108_),
    .B(_13255_),
    .X(_06000_));
 sky130_fd_sc_hd__nor2_4 _17039_ (.A(net340),
    .B(_06000_),
    .Y(\hash.CA1.S0.X[3] ));
 sky130_fd_sc_hd__inv_1 _17040_ (.A(_00658_),
    .Y(\hash.CA1.S0.X[0] ));
 sky130_fd_sc_hd__or3_4 _17041_ (.A(_13241_),
    .B(_05998_),
    .C(\hash.CA1.S0.X[0] ),
    .X(_06001_));
 sky130_fd_sc_hd__xor2_1 _17042_ (.A(\hash.CA1.S0.X[3] ),
    .B(_06001_),
    .X(_00683_));
 sky130_fd_sc_hd__clkinv_16 _17043_ (.A(net340),
    .Y(_06002_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1204 ();
 sky130_fd_sc_hd__a21o_4 _17048_ (.A1(_13240_),
    .A2(_13248_),
    .B1(_13247_),
    .X(_06007_));
 sky130_fd_sc_hd__a21oi_1 _17049_ (.A1(_13255_),
    .A2(_06007_),
    .B1(_13254_),
    .Y(_06008_));
 sky130_fd_sc_hd__xnor2_1 _17050_ (.A(_13262_),
    .B(_06008_),
    .Y(_06009_));
 sky130_fd_sc_hd__and2_4 _17051_ (.A(_06002_),
    .B(_06009_),
    .X(_06010_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1203 ();
 sky130_fd_sc_hd__a211oi_2 _17053_ (.A1(_13544_),
    .A2(_12109_),
    .B1(_06000_),
    .C1(net340),
    .Y(_06011_));
 sky130_fd_sc_hd__xor2_1 _17054_ (.A(_06010_),
    .B(_06011_),
    .X(_00684_));
 sky130_fd_sc_hd__nor2b_4 _17055_ (.A(_12108_),
    .B_N(_13255_),
    .Y(_06012_));
 sky130_fd_sc_hd__o21a_1 _17056_ (.A1(_13254_),
    .A2(_06012_),
    .B1(_13262_),
    .X(_06013_));
 sky130_fd_sc_hd__o21ai_2 _17057_ (.A1(_13261_),
    .A2(_06013_),
    .B1(_13269_),
    .Y(_06014_));
 sky130_fd_sc_hd__or3_4 _17058_ (.A(_13269_),
    .B(_13261_),
    .C(_06013_),
    .X(_06015_));
 sky130_fd_sc_hd__a21oi_4 _17059_ (.A1(_06014_),
    .A2(_06015_),
    .B1(net341),
    .Y(_06016_));
 sky130_fd_sc_hd__inv_2 _17060_ (.A(_06016_),
    .Y(\hash.CA1.S0.X[5] ));
 sky130_fd_sc_hd__nand4_1 _17061_ (.A(_06002_),
    .B(\hash.CA1.S0.X[3] ),
    .C(_06001_),
    .D(_06009_),
    .Y(_06017_));
 sky130_fd_sc_hd__xnor2_1 _17062_ (.A(_06016_),
    .B(_06017_),
    .Y(_00685_));
 sky130_fd_sc_hd__nor2_1 _17063_ (.A(net341),
    .B(_13276_),
    .Y(_06018_));
 sky130_fd_sc_hd__nor2b_1 _17064_ (.A(net341),
    .B_N(_13276_),
    .Y(_06019_));
 sky130_fd_sc_hd__or2_4 _17065_ (.A(_13254_),
    .B(_13261_),
    .X(_06020_));
 sky130_fd_sc_hd__a21oi_2 _17066_ (.A1(_13255_),
    .A2(_06007_),
    .B1(_06020_),
    .Y(_06021_));
 sky130_fd_sc_hd__o21ai_2 _17067_ (.A1(_13262_),
    .A2(_13261_),
    .B1(_13269_),
    .Y(_06022_));
 sky130_fd_sc_hd__o21bai_1 _17068_ (.A1(_06021_),
    .A2(_06022_),
    .B1_N(_13268_),
    .Y(_06023_));
 sky130_fd_sc_hd__mux2_8 _17069_ (.A0(_06018_),
    .A1(_06019_),
    .S(_06023_),
    .X(_06024_));
 sky130_fd_sc_hd__inv_4 _17070_ (.A(_06024_),
    .Y(\hash.CA1.S0.X[6] ));
 sky130_fd_sc_hd__nand3_2 _17071_ (.A(_06002_),
    .B(_06009_),
    .C(_06011_),
    .Y(_06025_));
 sky130_fd_sc_hd__nand2_1 _17072_ (.A(_06016_),
    .B(_06025_),
    .Y(_06026_));
 sky130_fd_sc_hd__xnor2_1 _17073_ (.A(\hash.CA1.S0.X[6] ),
    .B(_06026_),
    .Y(_00686_));
 sky130_fd_sc_hd__o21a_1 _17074_ (.A1(_13262_),
    .A2(_13261_),
    .B1(_13269_),
    .X(_06027_));
 sky130_fd_sc_hd__o211a_4 _17075_ (.A1(_06012_),
    .A2(_06020_),
    .B1(_06027_),
    .C1(_13276_),
    .X(_06028_));
 sky130_fd_sc_hd__a21o_4 _17076_ (.A1(_13276_),
    .A2(_13268_),
    .B1(_13275_),
    .X(_06029_));
 sky130_fd_sc_hd__or3_4 _17077_ (.A(_13283_),
    .B(_06028_),
    .C(_06029_),
    .X(_06030_));
 sky130_fd_sc_hd__o21ai_2 _17078_ (.A1(_06028_),
    .A2(_06029_),
    .B1(_13283_),
    .Y(_06031_));
 sky130_fd_sc_hd__nand3_4 _17079_ (.A(_06002_),
    .B(_06030_),
    .C(_06031_),
    .Y(_06032_));
 sky130_fd_sc_hd__inv_4 _17080_ (.A(_06032_),
    .Y(\hash.CA1.S0.X[7] ));
 sky130_fd_sc_hd__a31oi_2 _17081_ (.A1(_06016_),
    .A2(_06017_),
    .A3(_06024_),
    .B1(_06032_),
    .Y(_06033_));
 sky130_fd_sc_hd__nand3_1 _17082_ (.A(_06016_),
    .B(_06017_),
    .C(_06024_),
    .Y(_06034_));
 sky130_fd_sc_hd__nor2_1 _17083_ (.A(\hash.CA1.S0.X[7] ),
    .B(_06034_),
    .Y(_06035_));
 sky130_fd_sc_hd__nor2_1 _17084_ (.A(_06033_),
    .B(_06035_),
    .Y(_00687_));
 sky130_fd_sc_hd__nor2_1 _17085_ (.A(net341),
    .B(_13290_),
    .Y(_06036_));
 sky130_fd_sc_hd__nor2b_1 _17086_ (.A(net341),
    .B_N(_13290_),
    .Y(_06037_));
 sky130_fd_sc_hd__nor2_1 _17087_ (.A(_13268_),
    .B(_13275_),
    .Y(_06038_));
 sky130_fd_sc_hd__o21ai_0 _17088_ (.A1(_06021_),
    .A2(_06022_),
    .B1(_06038_),
    .Y(_06039_));
 sky130_fd_sc_hd__nor2_1 _17089_ (.A(_13276_),
    .B(_13275_),
    .Y(_06040_));
 sky130_fd_sc_hd__inv_1 _17090_ (.A(_06040_),
    .Y(_06041_));
 sky130_fd_sc_hd__a31oi_1 _17091_ (.A1(_13283_),
    .A2(_06039_),
    .A3(_06041_),
    .B1(_13282_),
    .Y(_06042_));
 sky130_fd_sc_hd__mux2_8 _17092_ (.A0(_06036_),
    .A1(_06037_),
    .S(_06042_),
    .X(_06043_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1202 ();
 sky130_fd_sc_hd__a31oi_2 _17094_ (.A1(_06016_),
    .A2(_06024_),
    .A3(_06025_),
    .B1(_06032_),
    .Y(_06044_));
 sky130_fd_sc_hd__xor2_1 _17095_ (.A(_06043_),
    .B(_06044_),
    .X(_00688_));
 sky130_fd_sc_hd__o211ai_1 _17096_ (.A1(_06012_),
    .A2(_06020_),
    .B1(_06027_),
    .C1(_13276_),
    .Y(_06045_));
 sky130_fd_sc_hd__nor3_4 _17097_ (.A(_13282_),
    .B(_13289_),
    .C(_06029_),
    .Y(_06046_));
 sky130_fd_sc_hd__o21a_4 _17098_ (.A1(_13283_),
    .A2(_13282_),
    .B1(_13290_),
    .X(_06047_));
 sky130_fd_sc_hd__nor2_1 _17099_ (.A(_13289_),
    .B(_06047_),
    .Y(_06048_));
 sky130_fd_sc_hd__a21oi_2 _17100_ (.A1(net1108),
    .A2(_06046_),
    .B1(_06048_),
    .Y(_06049_));
 sky130_fd_sc_hd__xnor2_2 _17101_ (.A(_13297_),
    .B(_06049_),
    .Y(_06050_));
 sky130_fd_sc_hd__nand2_8 _17102_ (.A(_06002_),
    .B(_06050_),
    .Y(\hash.CA1.S0.X[9] ));
 sky130_fd_sc_hd__nand2_1 _17103_ (.A(_06033_),
    .B(_06043_),
    .Y(_06051_));
 sky130_fd_sc_hd__xor2_1 _17104_ (.A(\hash.CA1.S0.X[9] ),
    .B(_06051_),
    .X(_00689_));
 sky130_fd_sc_hd__a21oi_2 _17105_ (.A1(_13297_),
    .A2(_13289_),
    .B1(_13282_),
    .Y(_06052_));
 sky130_fd_sc_hd__and2_0 _17106_ (.A(_06038_),
    .B(_06052_),
    .X(_06053_));
 sky130_fd_sc_hd__o21ai_2 _17107_ (.A1(_06021_),
    .A2(_06022_),
    .B1(_06053_),
    .Y(_06054_));
 sky130_fd_sc_hd__o21ai_4 _17108_ (.A1(_13289_),
    .A2(_06047_),
    .B1(_13297_),
    .Y(_06055_));
 sky130_fd_sc_hd__a21oi_2 _17109_ (.A1(_06040_),
    .A2(_06052_),
    .B1(_06055_),
    .Y(_06056_));
 sky130_fd_sc_hd__a21oi_2 _17110_ (.A1(_06054_),
    .A2(_06056_),
    .B1(_13296_),
    .Y(_06057_));
 sky130_fd_sc_hd__xnor2_4 _17111_ (.A(_13304_),
    .B(_06057_),
    .Y(_06058_));
 sky130_fd_sc_hd__nor2_4 _17112_ (.A(net340),
    .B(_06058_),
    .Y(_06059_));
 sky130_fd_sc_hd__inv_6 _17113_ (.A(_06059_),
    .Y(\hash.CA1.S0.X[10] ));
 sky130_fd_sc_hd__a21oi_1 _17114_ (.A1(_06043_),
    .A2(_06044_),
    .B1(\hash.CA1.S0.X[9] ),
    .Y(_06060_));
 sky130_fd_sc_hd__xnor2_1 _17115_ (.A(_06059_),
    .B(_06060_),
    .Y(_00659_));
 sky130_fd_sc_hd__inv_1 _17116_ (.A(_13304_),
    .Y(_06061_));
 sky130_fd_sc_hd__a211oi_4 _17117_ (.A1(_06046_),
    .A2(_06045_),
    .B1(_06061_),
    .C1(_06055_),
    .Y(_06062_));
 sky130_fd_sc_hd__a21o_1 _17118_ (.A1(_13304_),
    .A2(_13296_),
    .B1(_13303_),
    .X(_06063_));
 sky130_fd_sc_hd__nor2_1 _17119_ (.A(_06062_),
    .B(_06063_),
    .Y(_06064_));
 sky130_fd_sc_hd__xnor2_2 _17120_ (.A(_13311_),
    .B(_06064_),
    .Y(_06065_));
 sky130_fd_sc_hd__nand2_8 _17121_ (.A(_06002_),
    .B(_06065_),
    .Y(_06066_));
 sky130_fd_sc_hd__inv_1 _17122_ (.A(_06066_),
    .Y(\hash.CA1.S0.X[11] ));
 sky130_fd_sc_hd__a2111oi_2 _17123_ (.A1(_06033_),
    .A2(_06043_),
    .B1(\hash.CA1.S0.X[9] ),
    .C1(_06058_),
    .D1(net340),
    .Y(_06067_));
 sky130_fd_sc_hd__xor2_1 _17124_ (.A(_06066_),
    .B(_06067_),
    .X(_00660_));
 sky130_fd_sc_hd__or2_4 _17125_ (.A(_13311_),
    .B(_13310_),
    .X(_06068_));
 sky130_fd_sc_hd__o31ai_2 _17126_ (.A1(_13304_),
    .A2(_13303_),
    .A3(_13310_),
    .B1(_06068_),
    .Y(_06069_));
 sky130_fd_sc_hd__or3_1 _17127_ (.A(_13296_),
    .B(_13303_),
    .C(_13310_),
    .X(_06070_));
 sky130_fd_sc_hd__a21oi_2 _17128_ (.A1(_06056_),
    .A2(_06054_),
    .B1(_06070_),
    .Y(_06071_));
 sky130_fd_sc_hd__or2_4 _17129_ (.A(_06069_),
    .B(_06071_),
    .X(_06072_));
 sky130_fd_sc_hd__xor2_4 _17130_ (.A(_13318_),
    .B(_06072_),
    .X(_06073_));
 sky130_fd_sc_hd__nor2_4 _17131_ (.A(net340),
    .B(_06073_),
    .Y(\hash.CA1.S0.X[12] ));
 sky130_fd_sc_hd__a2111oi_0 _17132_ (.A1(_06043_),
    .A2(_06044_),
    .B1(\hash.CA1.S0.X[9] ),
    .C1(_06058_),
    .D1(net340),
    .Y(_06074_));
 sky130_fd_sc_hd__nor2_2 _17133_ (.A(_06066_),
    .B(_06074_),
    .Y(_06075_));
 sky130_fd_sc_hd__xor2_1 _17134_ (.A(\hash.CA1.S0.X[12] ),
    .B(_06075_),
    .X(_00661_));
 sky130_fd_sc_hd__or3_4 _17135_ (.A(_13310_),
    .B(_13317_),
    .C(_06063_),
    .X(_06076_));
 sky130_fd_sc_hd__a21o_1 _17136_ (.A1(_13318_),
    .A2(_06068_),
    .B1(_13317_),
    .X(_06077_));
 sky130_fd_sc_hd__o21ai_4 _17137_ (.A1(_06062_),
    .A2(_06076_),
    .B1(_06077_),
    .Y(_06078_));
 sky130_fd_sc_hd__xnor2_4 _17138_ (.A(_13325_),
    .B(_06078_),
    .Y(_06079_));
 sky130_fd_sc_hd__nor2_2 _17139_ (.A(net340),
    .B(_06079_),
    .Y(_06080_));
 sky130_fd_sc_hd__clkinv_1 _17140_ (.A(_06080_),
    .Y(\hash.CA1.S0.X[13] ));
 sky130_fd_sc_hd__nor4_2 _17141_ (.A(net340),
    .B(_06066_),
    .C(_06067_),
    .D(_06073_),
    .Y(_06081_));
 sky130_fd_sc_hd__xnor2_1 _17142_ (.A(\hash.CA1.S0.X[13] ),
    .B(_06081_),
    .Y(_00662_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1201 ();
 sky130_fd_sc_hd__clkinv_1 _17144_ (.A(_13332_),
    .Y(_06083_));
 sky130_fd_sc_hd__nor3_1 _17145_ (.A(_06083_),
    .B(_13317_),
    .C(_13324_),
    .Y(_06084_));
 sky130_fd_sc_hd__o21ai_0 _17146_ (.A1(_13318_),
    .A2(_13317_),
    .B1(_13325_),
    .Y(_06085_));
 sky130_fd_sc_hd__nand2b_1 _17147_ (.A_N(_13324_),
    .B(_06085_),
    .Y(_06086_));
 sky130_fd_sc_hd__nand2_1 _17148_ (.A(_13332_),
    .B(_06086_),
    .Y(_06087_));
 sky130_fd_sc_hd__nand2_1 _17149_ (.A(_13318_),
    .B(_13325_),
    .Y(_06088_));
 sky130_fd_sc_hd__a21oi_1 _17150_ (.A1(_13325_),
    .A2(_13317_),
    .B1(_13324_),
    .Y(_06089_));
 sky130_fd_sc_hd__o311ai_0 _17151_ (.A1(_06069_),
    .A2(_06071_),
    .A3(_06088_),
    .B1(_06089_),
    .C1(_06083_),
    .Y(_06090_));
 sky130_fd_sc_hd__a22oi_2 _17152_ (.A1(_06072_),
    .A2(_06084_),
    .B1(_06087_),
    .B2(_06090_),
    .Y(_06091_));
 sky130_fd_sc_hd__nand2_4 _17153_ (.A(_06002_),
    .B(_06091_),
    .Y(\hash.CA1.S0.X[14] ));
 sky130_fd_sc_hd__nand2_1 _17154_ (.A(\hash.CA1.S0.X[12] ),
    .B(_06075_),
    .Y(_06092_));
 sky130_fd_sc_hd__nand2_1 _17155_ (.A(_06080_),
    .B(_06092_),
    .Y(_06093_));
 sky130_fd_sc_hd__xnor2_1 _17156_ (.A(\hash.CA1.S0.X[14] ),
    .B(_06093_),
    .Y(_00663_));
 sky130_fd_sc_hd__a21oi_2 _17157_ (.A1(_13332_),
    .A2(_13324_),
    .B1(_13331_),
    .Y(_06094_));
 sky130_fd_sc_hd__nor2_1 _17158_ (.A(_13325_),
    .B(_13324_),
    .Y(_06095_));
 sky130_fd_sc_hd__nor2_1 _17159_ (.A(_06083_),
    .B(_06095_),
    .Y(_06096_));
 sky130_fd_sc_hd__nor2_1 _17160_ (.A(_13331_),
    .B(_06096_),
    .Y(_06097_));
 sky130_fd_sc_hd__a21oi_2 _17161_ (.A1(_06078_),
    .A2(_06094_),
    .B1(_06097_),
    .Y(_06098_));
 sky130_fd_sc_hd__xnor2_4 _17162_ (.A(_13339_),
    .B(_06098_),
    .Y(_06099_));
 sky130_fd_sc_hd__nand2_8 _17163_ (.A(_06002_),
    .B(_06099_),
    .Y(\hash.CA1.S0.X[15] ));
 sky130_fd_sc_hd__or3_1 _17164_ (.A(\hash.CA1.S0.X[13] ),
    .B(_06081_),
    .C(\hash.CA1.S0.X[14] ),
    .X(_06100_));
 sky130_fd_sc_hd__xnor2_1 _17165_ (.A(\hash.CA1.S0.X[15] ),
    .B(_06100_),
    .Y(_00664_));
 sky130_fd_sc_hd__or4_4 _17166_ (.A(_06083_),
    .B(_06069_),
    .C(_06088_),
    .D(_06071_),
    .X(_06101_));
 sky130_fd_sc_hd__a21o_4 _17167_ (.A1(_13325_),
    .A2(_13317_),
    .B1(_13324_),
    .X(_06102_));
 sky130_fd_sc_hd__nand2_2 _17168_ (.A(_13332_),
    .B(_06102_),
    .Y(_06103_));
 sky130_fd_sc_hd__nor2_1 _17169_ (.A(_13331_),
    .B(_13338_),
    .Y(_06104_));
 sky130_fd_sc_hd__nor2_1 _17170_ (.A(_13339_),
    .B(_13338_),
    .Y(_06105_));
 sky130_fd_sc_hd__a31oi_4 _17171_ (.A1(_06101_),
    .A2(_06103_),
    .A3(_06104_),
    .B1(_06105_),
    .Y(_06106_));
 sky130_fd_sc_hd__xor2_4 _17172_ (.A(_13346_),
    .B(_06106_),
    .X(_06107_));
 sky130_fd_sc_hd__nor2_4 _17173_ (.A(net340),
    .B(_06107_),
    .Y(_06108_));
 sky130_fd_sc_hd__inv_4 _17174_ (.A(_06108_),
    .Y(\hash.CA1.S0.X[16] ));
 sky130_fd_sc_hd__nand4_1 _17175_ (.A(_06002_),
    .B(_06080_),
    .C(_06091_),
    .D(_06099_),
    .Y(_06109_));
 sky130_fd_sc_hd__a21oi_2 _17176_ (.A1(\hash.CA1.S0.X[12] ),
    .A2(_06075_),
    .B1(_06109_),
    .Y(_06110_));
 sky130_fd_sc_hd__xnor2_1 _17177_ (.A(_06108_),
    .B(_06110_),
    .Y(_00665_));
 sky130_fd_sc_hd__inv_1 _17178_ (.A(_13345_),
    .Y(_06111_));
 sky130_fd_sc_hd__o21ai_2 _17179_ (.A1(_13331_),
    .A2(_06096_),
    .B1(_13339_),
    .Y(_06112_));
 sky130_fd_sc_hd__a21oi_1 _17180_ (.A1(_06078_),
    .A2(_06094_),
    .B1(_06112_),
    .Y(_06113_));
 sky130_fd_sc_hd__o21ai_1 _17181_ (.A1(_13338_),
    .A2(_06113_),
    .B1(_13346_),
    .Y(_06114_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1200 ();
 sky130_fd_sc_hd__a21boi_2 _17183_ (.A1(_06111_),
    .A2(_06114_),
    .B1_N(_13353_),
    .Y(_06116_));
 sky130_fd_sc_hd__nor3b_2 _17184_ (.A(_13353_),
    .B(_13345_),
    .C_N(_06114_),
    .Y(_06117_));
 sky130_fd_sc_hd__nor3_4 _17185_ (.A(net346),
    .B(_06116_),
    .C(_06117_),
    .Y(\hash.CA1.S0.X[17] ));
 sky130_fd_sc_hd__or3_4 _17186_ (.A(_06081_),
    .B(_06107_),
    .C(_06109_),
    .X(_06118_));
 sky130_fd_sc_hd__xor2_1 _17187_ (.A(\hash.CA1.S0.X[17] ),
    .B(_06118_),
    .X(_00666_));
 sky130_fd_sc_hd__a21o_1 _17188_ (.A1(_13353_),
    .A2(_13345_),
    .B1(_13352_),
    .X(_06119_));
 sky130_fd_sc_hd__a31oi_1 _17189_ (.A1(_13346_),
    .A2(_13353_),
    .A3(_06106_),
    .B1(_06119_),
    .Y(_06120_));
 sky130_fd_sc_hd__xnor2_2 _17190_ (.A(_13360_),
    .B(_06120_),
    .Y(_06121_));
 sky130_fd_sc_hd__nand2_4 _17191_ (.A(_06002_),
    .B(_06121_),
    .Y(_06122_));
 sky130_fd_sc_hd__inv_6 _17192_ (.A(_06122_),
    .Y(\hash.CA1.S0.X[18] ));
 sky130_fd_sc_hd__nand2_4 _17193_ (.A(_06108_),
    .B(_06110_),
    .Y(_06123_));
 sky130_fd_sc_hd__nand2_1 _17194_ (.A(\hash.CA1.S0.X[17] ),
    .B(_06123_),
    .Y(_06124_));
 sky130_fd_sc_hd__xnor2_1 _17195_ (.A(\hash.CA1.S0.X[18] ),
    .B(_06124_),
    .Y(_00667_));
 sky130_fd_sc_hd__nand2_2 _17196_ (.A(_13346_),
    .B(_13353_),
    .Y(_06125_));
 sky130_fd_sc_hd__nand3_1 _17197_ (.A(_13339_),
    .B(_13346_),
    .C(_13353_),
    .Y(_06126_));
 sky130_fd_sc_hd__nand3_1 _17198_ (.A(_13346_),
    .B(_13353_),
    .C(_13338_),
    .Y(_06127_));
 sky130_fd_sc_hd__o21ai_2 _17199_ (.A1(_06094_),
    .A2(_06126_),
    .B1(_06127_),
    .Y(_06128_));
 sky130_fd_sc_hd__nor2_1 _17200_ (.A(_06119_),
    .B(_06128_),
    .Y(_06129_));
 sky130_fd_sc_hd__o31ai_1 _17201_ (.A1(_06078_),
    .A2(_06112_),
    .A3(_06125_),
    .B1(_06129_),
    .Y(_06130_));
 sky130_fd_sc_hd__a21oi_1 _17202_ (.A1(_13360_),
    .A2(_06130_),
    .B1(_13359_),
    .Y(_06131_));
 sky130_fd_sc_hd__xnor2_2 _17203_ (.A(_13367_),
    .B(_06131_),
    .Y(_06132_));
 sky130_fd_sc_hd__nor2_4 _17204_ (.A(net341),
    .B(_06132_),
    .Y(_06133_));
 sky130_fd_sc_hd__clkinvlp_2 _17205_ (.A(_06133_),
    .Y(\hash.CA1.S0.X[19] ));
 sky130_fd_sc_hd__nand2_1 _17206_ (.A(\hash.CA1.S0.X[17] ),
    .B(_06118_),
    .Y(_06134_));
 sky130_fd_sc_hd__o21ai_2 _17207_ (.A1(_06134_),
    .A2(_06122_),
    .B1(_06133_),
    .Y(_06135_));
 sky130_fd_sc_hd__or3_1 _17208_ (.A(_06134_),
    .B(_06122_),
    .C(_06133_),
    .X(_06136_));
 sky130_fd_sc_hd__nand2_1 _17209_ (.A(_06135_),
    .B(_06136_),
    .Y(_00668_));
 sky130_fd_sc_hd__a21oi_2 _17210_ (.A1(_13332_),
    .A2(_06102_),
    .B1(_13331_),
    .Y(_06137_));
 sky130_fd_sc_hd__nand2_1 _17211_ (.A(_13360_),
    .B(_13367_),
    .Y(_06138_));
 sky130_fd_sc_hd__nor2_1 _17212_ (.A(_06125_),
    .B(_06138_),
    .Y(_06139_));
 sky130_fd_sc_hd__nand2_2 _17213_ (.A(_13339_),
    .B(_06139_),
    .Y(_06140_));
 sky130_fd_sc_hd__a21oi_4 _17214_ (.A1(_06101_),
    .A2(_06137_),
    .B1(_06140_),
    .Y(_06141_));
 sky130_fd_sc_hd__a21oi_1 _17215_ (.A1(_13353_),
    .A2(_13345_),
    .B1(_13352_),
    .Y(_06142_));
 sky130_fd_sc_hd__a21boi_0 _17216_ (.A1(_06142_),
    .A2(_06127_),
    .B1_N(_13360_),
    .Y(_06143_));
 sky130_fd_sc_hd__o21ai_2 _17217_ (.A1(_13359_),
    .A2(_06143_),
    .B1(_13367_),
    .Y(_06144_));
 sky130_fd_sc_hd__nand2b_4 _17218_ (.A_N(_13366_),
    .B(_06144_),
    .Y(_06145_));
 sky130_fd_sc_hd__or3_1 _17219_ (.A(_13374_),
    .B(_06141_),
    .C(_06145_),
    .X(_06146_));
 sky130_fd_sc_hd__o21ai_0 _17220_ (.A1(_06141_),
    .A2(_06145_),
    .B1(_13374_),
    .Y(_06147_));
 sky130_fd_sc_hd__and3_4 _17221_ (.A(_06002_),
    .B(_06146_),
    .C(_06147_),
    .X(_06148_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1199 ();
 sky130_fd_sc_hd__a31oi_2 _17223_ (.A1(\hash.CA1.S0.X[17] ),
    .A2(\hash.CA1.S0.X[18] ),
    .A3(_06123_),
    .B1(\hash.CA1.S0.X[19] ),
    .Y(_06149_));
 sky130_fd_sc_hd__xnor2_1 _17224_ (.A(_06148_),
    .B(_06149_),
    .Y(_00670_));
 sky130_fd_sc_hd__nor4_4 _17225_ (.A(_06128_),
    .B(_13366_),
    .C(_06119_),
    .D(_13359_),
    .Y(_06150_));
 sky130_fd_sc_hd__o31ai_4 _17226_ (.A1(_06078_),
    .A2(_06112_),
    .A3(_06125_),
    .B1(_06150_),
    .Y(_06151_));
 sky130_fd_sc_hd__o21ai_2 _17227_ (.A1(_13360_),
    .A2(_13359_),
    .B1(_13367_),
    .Y(_06152_));
 sky130_fd_sc_hd__nand2b_4 _17228_ (.A_N(_13366_),
    .B(_06152_),
    .Y(_06153_));
 sky130_fd_sc_hd__a31o_4 _17229_ (.A1(net1091),
    .A2(_13374_),
    .A3(_06153_),
    .B1(_13373_),
    .X(_06154_));
 sky130_fd_sc_hd__xor2_4 _17230_ (.A(_13381_),
    .B(_06154_),
    .X(_06155_));
 sky130_fd_sc_hd__and2_4 _17231_ (.A(_06002_),
    .B(_06155_),
    .X(_06156_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1198 ();
 sky130_fd_sc_hd__nand2_1 _17233_ (.A(_06135_),
    .B(_06148_),
    .Y(_06157_));
 sky130_fd_sc_hd__xnor2_1 _17234_ (.A(_06156_),
    .B(_06157_),
    .Y(_00671_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1197 ();
 sky130_fd_sc_hd__or3_4 _17236_ (.A(_13373_),
    .B(_13380_),
    .C(_06145_),
    .X(_06159_));
 sky130_fd_sc_hd__nor3_1 _17237_ (.A(_13374_),
    .B(_13373_),
    .C(_13380_),
    .Y(_06160_));
 sky130_fd_sc_hd__nor2_1 _17238_ (.A(_13381_),
    .B(_13380_),
    .Y(_06161_));
 sky130_fd_sc_hd__nor2_1 _17239_ (.A(_06160_),
    .B(_06161_),
    .Y(_06162_));
 sky130_fd_sc_hd__o21ai_2 _17240_ (.A1(_06141_),
    .A2(_06159_),
    .B1(_06162_),
    .Y(_06163_));
 sky130_fd_sc_hd__xor2_4 _17241_ (.A(_13388_),
    .B(_06163_),
    .X(_06164_));
 sky130_fd_sc_hd__nor2_4 _17242_ (.A(net341),
    .B(net1127),
    .Y(\hash.CA1.S0.X[22] ));
 sky130_fd_sc_hd__nand4_1 _17243_ (.A(_06002_),
    .B(_06146_),
    .C(_06147_),
    .D(_06155_),
    .Y(_06165_));
 sky130_fd_sc_hd__nor2_1 _17244_ (.A(_06149_),
    .B(_06165_),
    .Y(_06166_));
 sky130_fd_sc_hd__xor2_1 _17245_ (.A(\hash.CA1.S0.X[22] ),
    .B(_06166_),
    .X(_00672_));
 sky130_fd_sc_hd__a21o_1 _17246_ (.A1(_13381_),
    .A2(_06154_),
    .B1(_13380_),
    .X(_06167_));
 sky130_fd_sc_hd__a211o_4 _17247_ (.A1(_13388_),
    .A2(_06167_),
    .B1(_13387_),
    .C1(_13395_),
    .X(_06168_));
 sky130_fd_sc_hd__a211o_4 _17248_ (.A1(_06154_),
    .A2(_13381_),
    .B1(_13387_),
    .C1(_13380_),
    .X(_06169_));
 sky130_fd_sc_hd__o21a_4 _17249_ (.A1(_13388_),
    .A2(_13387_),
    .B1(_13395_),
    .X(_06170_));
 sky130_fd_sc_hd__a21oi_2 _17250_ (.A1(_06169_),
    .A2(_06170_),
    .B1(net341),
    .Y(_06171_));
 sky130_fd_sc_hd__nand2_8 _17251_ (.A(_06168_),
    .B(_06171_),
    .Y(_06172_));
 sky130_fd_sc_hd__inv_2 _17252_ (.A(_06172_),
    .Y(\hash.CA1.S0.X[23] ));
 sky130_fd_sc_hd__nor2_1 _17253_ (.A(net1127),
    .B(_06165_),
    .Y(_06173_));
 sky130_fd_sc_hd__nand2_1 _17254_ (.A(_06135_),
    .B(_06173_),
    .Y(_06174_));
 sky130_fd_sc_hd__xnor2_1 _17255_ (.A(\hash.CA1.S0.X[23] ),
    .B(_06174_),
    .Y(_00673_));
 sky130_fd_sc_hd__inv_1 _17256_ (.A(_13387_),
    .Y(_06175_));
 sky130_fd_sc_hd__o211ai_1 _17257_ (.A1(_06141_),
    .A2(_06159_),
    .B1(_06162_),
    .C1(_13388_),
    .Y(_06176_));
 sky130_fd_sc_hd__a21boi_2 _17258_ (.A1(_06175_),
    .A2(_06176_),
    .B1_N(_13395_),
    .Y(_06177_));
 sky130_fd_sc_hd__o21ai_1 _17259_ (.A1(_13394_),
    .A2(_06177_),
    .B1(_13402_),
    .Y(_06178_));
 sky130_fd_sc_hd__o311a_4 _17260_ (.A1(_13402_),
    .A2(_13394_),
    .A3(_06177_),
    .B1(_06178_),
    .C1(_06002_),
    .X(_06179_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1196 ();
 sky130_fd_sc_hd__nor4_2 _17262_ (.A(_06149_),
    .B(net1127),
    .C(_06165_),
    .D(_06172_),
    .Y(_06180_));
 sky130_fd_sc_hd__xor2_1 _17263_ (.A(_06179_),
    .B(_06180_),
    .X(_00674_));
 sky130_fd_sc_hd__clkinv_1 _17264_ (.A(_13409_),
    .Y(_06181_));
 sky130_fd_sc_hd__a2111o_2 _17265_ (.A1(_06169_),
    .A2(_06170_),
    .B1(_06181_),
    .C1(_13394_),
    .D1(_13401_),
    .X(_06182_));
 sky130_fd_sc_hd__inv_1 _17266_ (.A(_13402_),
    .Y(_06183_));
 sky130_fd_sc_hd__nor2_2 _17267_ (.A(_06183_),
    .B(_13409_),
    .Y(_06184_));
 sky130_fd_sc_hd__nand3_2 _17268_ (.A(_06169_),
    .B(_06170_),
    .C(_06184_),
    .Y(_06185_));
 sky130_fd_sc_hd__nor3_1 _17269_ (.A(_13402_),
    .B(_06181_),
    .C(_13401_),
    .Y(_06186_));
 sky130_fd_sc_hd__a221oi_2 _17270_ (.A1(_06181_),
    .A2(_13401_),
    .B1(_06184_),
    .B2(_13394_),
    .C1(_06186_),
    .Y(_06187_));
 sky130_fd_sc_hd__nand4_1 _17271_ (.A(_06002_),
    .B(_06182_),
    .C(_06185_),
    .D(_06187_),
    .Y(\hash.CA1.S0.X[25] ));
 sky130_fd_sc_hd__and4_4 _17272_ (.A(_06135_),
    .B(\hash.CA1.S0.X[23] ),
    .C(_06173_),
    .D(_06179_),
    .X(_06188_));
 sky130_fd_sc_hd__xnor2_1 _17273_ (.A(net1049),
    .B(_06188_),
    .Y(_00675_));
 sky130_fd_sc_hd__nand3_1 _17274_ (.A(_13388_),
    .B(_13395_),
    .C(_13402_),
    .Y(_06189_));
 sky130_fd_sc_hd__nand2_1 _17275_ (.A(_13381_),
    .B(_13409_),
    .Y(_06190_));
 sky130_fd_sc_hd__nor2_2 _17276_ (.A(_06189_),
    .B(_06190_),
    .Y(_06191_));
 sky130_fd_sc_hd__o211a_4 _17277_ (.A1(_06141_),
    .A2(_06145_),
    .B1(_06191_),
    .C1(_13374_),
    .X(_06192_));
 sky130_fd_sc_hd__a21oi_1 _17278_ (.A1(_13395_),
    .A2(_13387_),
    .B1(_13394_),
    .Y(_06193_));
 sky130_fd_sc_hd__a41oi_1 _17279_ (.A1(_13388_),
    .A2(_13395_),
    .A3(_13402_),
    .A4(_13380_),
    .B1(_13401_),
    .Y(_06194_));
 sky130_fd_sc_hd__o21ai_0 _17280_ (.A1(_06183_),
    .A2(_06193_),
    .B1(_06194_),
    .Y(_06195_));
 sky130_fd_sc_hd__a21oi_1 _17281_ (.A1(_13409_),
    .A2(_06195_),
    .B1(_13408_),
    .Y(_06196_));
 sky130_fd_sc_hd__nand2_1 _17282_ (.A(_13373_),
    .B(_06191_),
    .Y(_06197_));
 sky130_fd_sc_hd__nand2_2 _17283_ (.A(_06196_),
    .B(_06197_),
    .Y(_06198_));
 sky130_fd_sc_hd__nor3_2 _17284_ (.A(_13416_),
    .B(_06192_),
    .C(_06198_),
    .Y(_06199_));
 sky130_fd_sc_hd__o21a_4 _17285_ (.A1(_06192_),
    .A2(_06198_),
    .B1(_13416_),
    .X(_06200_));
 sky130_fd_sc_hd__nor3_4 _17286_ (.A(net341),
    .B(_06199_),
    .C(_06200_),
    .Y(_06201_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1195 ();
 sky130_fd_sc_hd__a21oi_1 _17288_ (.A1(_06179_),
    .A2(_06180_),
    .B1(\hash.CA1.S0.X[25] ),
    .Y(_06202_));
 sky130_fd_sc_hd__xnor2_1 _17289_ (.A(_06201_),
    .B(_06202_),
    .Y(_00676_));
 sky130_fd_sc_hd__and3_1 _17290_ (.A(_13374_),
    .B(_13416_),
    .C(_06191_),
    .X(_06203_));
 sky130_fd_sc_hd__nand3_2 _17291_ (.A(_06153_),
    .B(_06151_),
    .C(_06203_),
    .Y(_06204_));
 sky130_fd_sc_hd__inv_1 _17292_ (.A(_13416_),
    .Y(_06205_));
 sky130_fd_sc_hd__nand3_1 _17293_ (.A(_13416_),
    .B(_13373_),
    .C(_06191_),
    .Y(_06206_));
 sky130_fd_sc_hd__o21ai_0 _17294_ (.A1(_06205_),
    .A2(_06196_),
    .B1(_06206_),
    .Y(_06207_));
 sky130_fd_sc_hd__inv_1 _17295_ (.A(_06207_),
    .Y(_06208_));
 sky130_fd_sc_hd__nand3b_1 _17296_ (.A_N(_13415_),
    .B(_06204_),
    .C(_06208_),
    .Y(_06209_));
 sky130_fd_sc_hd__xor2_1 _17297_ (.A(_13423_),
    .B(_06209_),
    .X(_06210_));
 sky130_fd_sc_hd__or2_4 _17298_ (.A(net341),
    .B(_06210_),
    .X(_06211_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1194 ();
 sky130_fd_sc_hd__nand3_4 _17300_ (.A(_06182_),
    .B(_06185_),
    .C(_06187_),
    .Y(_06212_));
 sky130_fd_sc_hd__o21ai_0 _17301_ (.A1(_06212_),
    .A2(_06188_),
    .B1(_06201_),
    .Y(_06213_));
 sky130_fd_sc_hd__xor2_1 _17302_ (.A(_06211_),
    .B(_06213_),
    .X(_00677_));
 sky130_fd_sc_hd__o21a_1 _17303_ (.A1(_13415_),
    .A2(_06200_),
    .B1(_13423_),
    .X(_06214_));
 sky130_fd_sc_hd__nor3_1 _17304_ (.A(_13430_),
    .B(_13422_),
    .C(_06214_),
    .Y(_06215_));
 sky130_fd_sc_hd__or2_4 _17305_ (.A(_13423_),
    .B(_13422_),
    .X(_06216_));
 sky130_fd_sc_hd__o311a_4 _17306_ (.A1(_13415_),
    .A2(_13422_),
    .A3(_06200_),
    .B1(_06216_),
    .C1(_13430_),
    .X(_06217_));
 sky130_fd_sc_hd__or3_4 _17307_ (.A(net341),
    .B(_06215_),
    .C(_06217_),
    .X(_06218_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1193 ();
 sky130_fd_sc_hd__a21o_1 _17309_ (.A1(_06212_),
    .A2(_06201_),
    .B1(_06211_),
    .X(_06220_));
 sky130_fd_sc_hd__a31o_4 _17310_ (.A1(_06179_),
    .A2(_06180_),
    .A3(_06201_),
    .B1(_06220_),
    .X(_06221_));
 sky130_fd_sc_hd__xnor2_1 _17311_ (.A(_06218_),
    .B(_06221_),
    .Y(_00678_));
 sky130_fd_sc_hd__nor3_1 _17312_ (.A(_13415_),
    .B(_13422_),
    .C(_13429_),
    .Y(_06222_));
 sky130_fd_sc_hd__a21oi_1 _17313_ (.A1(_13430_),
    .A2(_06216_),
    .B1(_13429_),
    .Y(_06223_));
 sky130_fd_sc_hd__a31oi_4 _17314_ (.A1(_06208_),
    .A2(_06204_),
    .A3(_06222_),
    .B1(_06223_),
    .Y(_06224_));
 sky130_fd_sc_hd__xor2_1 _17315_ (.A(_13437_),
    .B(_06224_),
    .X(_06225_));
 sky130_fd_sc_hd__nor2_4 _17316_ (.A(net341),
    .B(_06225_),
    .Y(_06226_));
 sky130_fd_sc_hd__inv_4 _17317_ (.A(_06226_),
    .Y(\hash.CA1.S0.X[29] ));
 sky130_fd_sc_hd__and3b_1 _17318_ (.A_N(_06172_),
    .B(_06173_),
    .C(_06201_),
    .X(_06227_));
 sky130_fd_sc_hd__nand3_1 _17319_ (.A(_06135_),
    .B(_06179_),
    .C(_06227_),
    .Y(_06228_));
 sky130_fd_sc_hd__a21oi_1 _17320_ (.A1(_06212_),
    .A2(_06201_),
    .B1(_06211_),
    .Y(_06229_));
 sky130_fd_sc_hd__a21oi_2 _17321_ (.A1(_06228_),
    .A2(_06229_),
    .B1(_06218_),
    .Y(_06230_));
 sky130_fd_sc_hd__xnor2_1 _17322_ (.A(\hash.CA1.S0.X[29] ),
    .B(_06230_),
    .Y(_00679_));
 sky130_fd_sc_hd__o21a_1 _17323_ (.A1(_13429_),
    .A2(_06217_),
    .B1(_13437_),
    .X(_06231_));
 sky130_fd_sc_hd__o21ai_2 _17324_ (.A1(_13436_),
    .A2(_06231_),
    .B1(_13444_),
    .Y(_06232_));
 sky130_fd_sc_hd__or3_4 _17325_ (.A(_13444_),
    .B(_13436_),
    .C(_06231_),
    .X(_06233_));
 sky130_fd_sc_hd__a21o_4 _17326_ (.A1(_06233_),
    .A2(_06232_),
    .B1(net341),
    .X(_06234_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1192 ();
 sky130_fd_sc_hd__inv_1 _17328_ (.A(_06218_),
    .Y(\hash.CA1.S0.X[28] ));
 sky130_fd_sc_hd__a21o_1 _17329_ (.A1(\hash.CA1.S0.X[28] ),
    .A2(_06221_),
    .B1(\hash.CA1.S0.X[29] ),
    .X(_06235_));
 sky130_fd_sc_hd__xnor2_1 _17330_ (.A(_06234_),
    .B(_06235_),
    .Y(_00681_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1191 ();
 sky130_fd_sc_hd__maj3_1 _17332_ (.A(\hash.CA2.b_dash[31] ),
    .B(\hash.CA2.a_dash[31] ),
    .C(net1078),
    .X(_06237_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1190 ();
 sky130_fd_sc_hd__mux2i_1 _17334_ (.A0(\hash.CA2.f_dash[31] ),
    .A1(\hash.CA2.e_dash[31] ),
    .S(\hash.CA2.S1.X[31] ),
    .Y(_06239_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1187 ();
 sky130_fd_sc_hd__xor2_1 _17338_ (.A(\hash.CA2.S1.X[5] ),
    .B(\hash.CA2.S1.X[24] ),
    .X(_06243_));
 sky130_fd_sc_hd__xnor2_1 _17339_ (.A(\hash.CA2.S1.X[10] ),
    .B(_06243_),
    .Y(_06244_));
 sky130_fd_sc_hd__xnor2_2 _17340_ (.A(_06239_),
    .B(_06244_),
    .Y(_06245_));
 sky130_fd_sc_hd__o211ai_1 _17341_ (.A1(_04723_),
    .A2(_04749_),
    .B1(_04775_),
    .C1(_04751_),
    .Y(_06246_));
 sky130_fd_sc_hd__a31o_4 _17342_ (.A1(_13441_),
    .A2(_04776_),
    .A3(_06246_),
    .B1(_13440_),
    .X(_06247_));
 sky130_fd_sc_hd__xor2_4 _17343_ (.A(_06245_),
    .B(_06247_),
    .X(_06248_));
 sky130_fd_sc_hd__and3_1 _17344_ (.A(_04457_),
    .B(_04461_),
    .C(_04590_),
    .X(_06249_));
 sky130_fd_sc_hd__a21boi_0 _17345_ (.A1(_04457_),
    .A2(_04461_),
    .B1_N(_04592_),
    .Y(_06250_));
 sky130_fd_sc_hd__inv_1 _17346_ (.A(_04595_),
    .Y(_06251_));
 sky130_fd_sc_hd__xnor2_1 _17347_ (.A(\hash.CA2.p4[31] ),
    .B(_12360_),
    .Y(_06252_));
 sky130_fd_sc_hd__xnor2_1 _17348_ (.A(_12082_),
    .B(_12356_),
    .Y(_06253_));
 sky130_fd_sc_hd__xnor2_1 _17349_ (.A(_06252_),
    .B(_06253_),
    .Y(_06254_));
 sky130_fd_sc_hd__xnor3_1 _17350_ (.A(_12948_),
    .B(net1096),
    .C(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__or4_4 _17351_ (.A(_06249_),
    .B(_06250_),
    .C(_06251_),
    .D(_06255_),
    .X(_06256_));
 sky130_fd_sc_hd__o31ai_1 _17352_ (.A1(_06249_),
    .A2(_06250_),
    .A3(_06251_),
    .B1(_06255_),
    .Y(_06257_));
 sky130_fd_sc_hd__nand2_2 _17353_ (.A(_06256_),
    .B(_06257_),
    .Y(_06258_));
 sky130_fd_sc_hd__nand2_1 _17354_ (.A(_13444_),
    .B(_13436_),
    .Y(_06259_));
 sky130_fd_sc_hd__inv_1 _17355_ (.A(_13443_),
    .Y(_06260_));
 sky130_fd_sc_hd__a22oi_1 _17356_ (.A1(_06256_),
    .A2(_06257_),
    .B1(_06259_),
    .B2(_06260_),
    .Y(_06261_));
 sky130_fd_sc_hd__a41o_1 _17357_ (.A1(_13437_),
    .A2(_13444_),
    .A3(_06224_),
    .A4(_06258_),
    .B1(_06261_),
    .X(_06262_));
 sky130_fd_sc_hd__nor4_1 _17358_ (.A(_13436_),
    .B(_13443_),
    .C(_06224_),
    .D(_06258_),
    .Y(_06263_));
 sky130_fd_sc_hd__nor4_1 _17359_ (.A(_13437_),
    .B(_13436_),
    .C(_13443_),
    .D(_06258_),
    .Y(_06264_));
 sky130_fd_sc_hd__nor3_1 _17360_ (.A(_13444_),
    .B(_13443_),
    .C(_06258_),
    .Y(_06265_));
 sky130_fd_sc_hd__or4_4 _17361_ (.A(_06262_),
    .B(_06263_),
    .C(_06264_),
    .D(_06265_),
    .X(_06266_));
 sky130_fd_sc_hd__xor2_2 _17362_ (.A(_06248_),
    .B(_06266_),
    .X(_06267_));
 sky130_fd_sc_hd__xnor2_2 _17363_ (.A(_06237_),
    .B(_06267_),
    .Y(_06268_));
 sky130_fd_sc_hd__nand2_8 _17364_ (.A(_06002_),
    .B(_06268_),
    .Y(_06269_));
 sky130_fd_sc_hd__inv_1 _17365_ (.A(_06269_),
    .Y(\hash.CA1.S0.X[31] ));
 sky130_fd_sc_hd__nor3_1 _17366_ (.A(\hash.CA1.S0.X[29] ),
    .B(_06230_),
    .C(_06234_),
    .Y(_06270_));
 sky130_fd_sc_hd__xor2_1 _17367_ (.A(_06269_),
    .B(_06270_),
    .X(_00682_));
 sky130_fd_sc_hd__xor2_1 _17368_ (.A(\hash.CA1.S0.X[3] ),
    .B(\hash.CA1.S0.X[14] ),
    .X(_06271_));
 sky130_fd_sc_hd__xnor2_1 _17369_ (.A(_06172_),
    .B(_06271_),
    .Y(_13548_));
 sky130_fd_sc_hd__inv_1 _17370_ (.A(_13548_),
    .Y(_12881_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1184 ();
 sky130_fd_sc_hd__nor2b_4 _17374_ (.A(net340),
    .B_N(_12082_),
    .Y(\hash.CA1.b[1] ));
 sky130_fd_sc_hd__a21oi_1 _17375_ (.A1(\hash.CA2.a_dash[1] ),
    .A2(_13241_),
    .B1(_12082_),
    .Y(_06275_));
 sky130_fd_sc_hd__nor2_1 _17376_ (.A(\hash.CA2.a_dash[1] ),
    .B(_13241_),
    .Y(_06276_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1183 ();
 sky130_fd_sc_hd__o21ai_0 _17378_ (.A1(_06275_),
    .A2(_06276_),
    .B1(_06002_),
    .Y(_13547_));
 sky130_fd_sc_hd__inv_1 _17379_ (.A(_13547_),
    .Y(_12880_));
 sky130_fd_sc_hd__nor2b_4 _17380_ (.A(net340),
    .B_N(\hash.CA2.a_dash[0] ),
    .Y(\hash.CA1.c[0] ));
 sky130_fd_sc_hd__nand2b_1 _17381_ (.A_N(_04421_),
    .B(_06002_),
    .Y(\hash.CA1.b[2] ));
 sky130_fd_sc_hd__nor2b_4 _17382_ (.A(net340),
    .B_N(\hash.CA2.a_dash[2] ),
    .Y(_13673_));
 sky130_fd_sc_hd__and2_0 _17383_ (.A(_06002_),
    .B(_04470_),
    .X(\hash.CA1.b[3] ));
 sky130_fd_sc_hd__nor2b_4 _17384_ (.A(net340),
    .B_N(\hash.CA2.a_dash[3] ),
    .Y(_13679_));
 sky130_fd_sc_hd__and2_4 _17385_ (.A(_06002_),
    .B(_04487_),
    .X(\hash.CA1.b[4] ));
 sky130_fd_sc_hd__and2_4 _17386_ (.A(_06002_),
    .B(_04501_),
    .X(\hash.CA1.b[5] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1182 ();
 sky130_fd_sc_hd__or2_4 _17388_ (.A(net341),
    .B(\hash.CA2.a_dash[5] ),
    .X(_13691_));
 sky130_fd_sc_hd__and2_4 _17389_ (.A(_06002_),
    .B(_04522_),
    .X(\hash.CA1.b[6] ));
 sky130_fd_sc_hd__or2_4 _17390_ (.A(net340),
    .B(\hash.CA2.a_dash[6] ),
    .X(_13697_));
 sky130_fd_sc_hd__nand2_2 _17391_ (.A(_06002_),
    .B(_04543_),
    .Y(\hash.CA1.b[7] ));
 sky130_fd_sc_hd__and2_4 _17392_ (.A(_06002_),
    .B(_04562_),
    .X(_06279_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1181 ();
 sky130_fd_sc_hd__or2_4 _17394_ (.A(net340),
    .B(_04580_),
    .X(_06280_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1180 ();
 sky130_fd_sc_hd__or2_4 _17396_ (.A(net340),
    .B(\hash.CA2.a_dash[9] ),
    .X(_13716_));
 sky130_fd_sc_hd__or2_4 _17397_ (.A(net341),
    .B(_04599_),
    .X(\hash.CA1.b[10] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1179 ();
 sky130_fd_sc_hd__nor2_4 _17399_ (.A(net340),
    .B(_04614_),
    .Y(_06282_));
 sky130_fd_sc_hd__inv_1 _17400_ (.A(_06282_),
    .Y(\hash.CA1.b[11] ));
 sky130_fd_sc_hd__and2_4 _17401_ (.A(_06002_),
    .B(_04623_),
    .X(_06283_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1178 ();
 sky130_fd_sc_hd__or2_0 _17403_ (.A(net341),
    .B(_04437_),
    .X(\hash.CA1.b[13] ));
 sky130_fd_sc_hd__or2_4 _17404_ (.A(net346),
    .B(\hash.CA2.a_dash[13] ),
    .X(_13740_));
 sky130_fd_sc_hd__nor2_1 _17405_ (.A(net341),
    .B(_04475_),
    .Y(\hash.CA1.b[14] ));
 sky130_fd_sc_hd__or2_4 _17406_ (.A(net341),
    .B(\hash.CA2.a_dash[14] ),
    .X(_13746_));
 sky130_fd_sc_hd__or2_4 _17407_ (.A(net341),
    .B(_04484_),
    .X(\hash.CA1.b[15] ));
 sky130_fd_sc_hd__or2_4 _17408_ (.A(net341),
    .B(\hash.CA2.a_dash[15] ),
    .X(_13753_));
 sky130_fd_sc_hd__nand2b_2 _17409_ (.A_N(_04503_),
    .B(_06002_),
    .Y(\hash.CA1.b[16] ));
 sky130_fd_sc_hd__or2_4 _17410_ (.A(net341),
    .B(_04520_),
    .X(\hash.CA1.b[17] ));
 sky130_fd_sc_hd__or2_4 _17411_ (.A(net341),
    .B(_04541_),
    .X(\hash.CA1.b[18] ));
 sky130_fd_sc_hd__and2_4 _17412_ (.A(_06002_),
    .B(_04559_),
    .X(_06284_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1177 ();
 sky130_fd_sc_hd__or2_4 _17414_ (.A(net341),
    .B(\hash.CA2.a_dash[19] ),
    .X(_13778_));
 sky130_fd_sc_hd__nor2_1 _17415_ (.A(net341),
    .B(_04681_),
    .Y(\hash.CA1.b[20] ));
 sky130_fd_sc_hd__nand4_1 _17416_ (.A(_06002_),
    .B(_04591_),
    .C(_04593_),
    .D(_04595_),
    .Y(\hash.CA1.b[21] ));
 sky130_fd_sc_hd__or2_4 _17417_ (.A(net343),
    .B(_04420_),
    .X(\hash.CA1.b[22] ));
 sky130_fd_sc_hd__and2_4 _17418_ (.A(_06002_),
    .B(_04467_),
    .X(_06285_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1176 ();
 sky130_fd_sc_hd__nand2_2 _17420_ (.A(_06002_),
    .B(_04481_),
    .Y(\hash.CA1.b[24] ));
 sky130_fd_sc_hd__nand2_4 _17421_ (.A(_06002_),
    .B(_04499_),
    .Y(\hash.CA1.b[25] ));
 sky130_fd_sc_hd__clkinv_1 _17422_ (.A(net1103),
    .Y(_06286_));
 sky130_fd_sc_hd__nor2_2 _17423_ (.A(net343),
    .B(_06286_),
    .Y(\hash.CA1.b[26] ));
 sky130_fd_sc_hd__or2_4 _17424_ (.A(net343),
    .B(\hash.CA2.a_dash[26] ),
    .X(_06287_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1175 ();
 sky130_fd_sc_hd__nor2_2 _17426_ (.A(net341),
    .B(net1069),
    .Y(_06288_));
 sky130_fd_sc_hd__inv_1 _17427_ (.A(_06288_),
    .Y(\hash.CA1.b[27] ));
 sky130_fd_sc_hd__or2_4 _17428_ (.A(net346),
    .B(\hash.CA2.a_dash[27] ),
    .X(_13827_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1174 ();
 sky130_fd_sc_hd__nand2_1 _17430_ (.A(_06002_),
    .B(_04662_),
    .Y(\hash.CA1.b[28] ));
 sky130_fd_sc_hd__or2_4 _17431_ (.A(net343),
    .B(\hash.CA2.a_dash[28] ),
    .X(_13834_));
 sky130_fd_sc_hd__or2_4 _17432_ (.A(net343),
    .B(\hash.CA2.a_dash[29] ),
    .X(_13840_));
 sky130_fd_sc_hd__nor2_1 _17433_ (.A(net341),
    .B(_04588_),
    .Y(\hash.CA1.b[30] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1173 ();
 sky130_fd_sc_hd__o21ai_0 _17435_ (.A1(_04608_),
    .A2(_04611_),
    .B1(_06002_),
    .Y(\hash.CA1.b[31] ));
 sky130_fd_sc_hd__nor2_4 _17436_ (.A(net344),
    .B(\hash.CA2.e_dash[1] ),
    .Y(_12368_));
 sky130_fd_sc_hd__nor2b_4 _17437_ (.A(net343),
    .B_N(\hash.CA2.e_dash[2] ),
    .Y(_12375_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1172 ();
 sky130_fd_sc_hd__nor2_4 _17439_ (.A(net343),
    .B(\hash.CA2.e_dash[3] ),
    .Y(_12383_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1171 ();
 sky130_fd_sc_hd__nor2b_4 _17441_ (.A(net343),
    .B_N(\hash.CA2.e_dash[4] ),
    .Y(_12386_));
 sky130_fd_sc_hd__nor2_4 _17442_ (.A(net343),
    .B(\hash.CA2.e_dash[5] ),
    .Y(_12391_));
 sky130_fd_sc_hd__nor2b_4 _17443_ (.A(net343),
    .B_N(\hash.CA2.e_dash[6] ),
    .Y(_12394_));
 sky130_fd_sc_hd__nor2_4 _17444_ (.A(net343),
    .B(\hash.CA2.e_dash[7] ),
    .Y(_12399_));
 sky130_fd_sc_hd__nor2_4 _17445_ (.A(net343),
    .B(\hash.CA2.e_dash[8] ),
    .Y(_12404_));
 sky130_fd_sc_hd__nor2b_4 _17446_ (.A(net343),
    .B_N(\hash.CA2.e_dash[9] ),
    .Y(_12407_));
 sky130_fd_sc_hd__nor2b_4 _17447_ (.A(net343),
    .B_N(\hash.CA2.e_dash[10] ),
    .Y(_12410_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1170 ();
 sky130_fd_sc_hd__nor2_4 _17449_ (.A(net346),
    .B(\hash.CA2.e_dash[11] ),
    .Y(_12415_));
 sky130_fd_sc_hd__nor2_4 _17450_ (.A(net346),
    .B(\hash.CA2.e_dash[12] ),
    .Y(_12420_));
 sky130_fd_sc_hd__nor2b_4 _17451_ (.A(net343),
    .B_N(\hash.CA2.e_dash[13] ),
    .Y(_12423_));
 sky130_fd_sc_hd__nor2_4 _17452_ (.A(net343),
    .B(\hash.CA2.e_dash[14] ),
    .Y(_12428_));
 sky130_fd_sc_hd__nor2_4 _17453_ (.A(net343),
    .B(\hash.CA2.e_dash[15] ),
    .Y(_12433_));
 sky130_fd_sc_hd__nor2_4 _17454_ (.A(net343),
    .B(\hash.CA2.e_dash[16] ),
    .Y(_12438_));
 sky130_fd_sc_hd__nor2_4 _17455_ (.A(net343),
    .B(\hash.CA2.e_dash[17] ),
    .Y(_12443_));
 sky130_fd_sc_hd__nor2b_4 _17456_ (.A(net343),
    .B_N(\hash.CA2.e_dash[18] ),
    .Y(_12446_));
 sky130_fd_sc_hd__clkinv_1 _17457_ (.A(\hash.CA2.e_dash[19] ),
    .Y(_06294_));
 sky130_fd_sc_hd__nor2_4 _17458_ (.A(net343),
    .B(_06294_),
    .Y(_12449_));
 sky130_fd_sc_hd__nor2b_4 _17459_ (.A(net342),
    .B_N(\hash.CA2.e_dash[20] ),
    .Y(_12452_));
 sky130_fd_sc_hd__nor2b_4 _17460_ (.A(net342),
    .B_N(\hash.CA2.e_dash[21] ),
    .Y(_12455_));
 sky130_fd_sc_hd__nor2b_4 _17461_ (.A(\hash.reset ),
    .B_N(\hash.CA2.e_dash[22] ),
    .Y(_12458_));
 sky130_fd_sc_hd__nor2_4 _17462_ (.A(net344),
    .B(\hash.CA2.e_dash[23] ),
    .Y(_12463_));
 sky130_fd_sc_hd__nor2_1 _17463_ (.A(net346),
    .B(\hash.CA2.e_dash[24] ),
    .Y(_12468_));
 sky130_fd_sc_hd__nor2_4 _17464_ (.A(net346),
    .B(\hash.CA2.e_dash[25] ),
    .Y(_12473_));
 sky130_fd_sc_hd__nor2_4 _17465_ (.A(net346),
    .B(\hash.CA2.e_dash[26] ),
    .Y(_12478_));
 sky130_fd_sc_hd__nor2_4 _17466_ (.A(net346),
    .B(\hash.CA2.e_dash[27] ),
    .Y(_12483_));
 sky130_fd_sc_hd__nor2_2 _17467_ (.A(net346),
    .B(\hash.CA2.e_dash[28] ),
    .Y(_12488_));
 sky130_fd_sc_hd__nor2b_4 _17468_ (.A(net345),
    .B_N(\hash.CA2.e_dash[29] ),
    .Y(_12491_));
 sky130_fd_sc_hd__nor2b_1 _17469_ (.A(net346),
    .B_N(\hash.CA2.e_dash[30] ),
    .Y(_12494_));
 sky130_fd_sc_hd__nor2b_4 _17470_ (.A(net343),
    .B_N(\hash.CA2.f_dash[1] ),
    .Y(_12505_));
 sky130_fd_sc_hd__nand2_8 _17471_ (.A(_06002_),
    .B(\hash.CA2.f_dash[2] ),
    .Y(_12667_));
 sky130_fd_sc_hd__inv_6 _17472_ (.A(_12667_),
    .Y(_12510_));
 sky130_fd_sc_hd__xor2_1 _17473_ (.A(_13848_),
    .B(_12510_),
    .X(_00896_));
 sky130_fd_sc_hd__nor2_4 _17474_ (.A(net344),
    .B(\hash.CA2.f_dash[3] ),
    .Y(_12515_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1169 ();
 sky130_fd_sc_hd__nand3_2 _17476_ (.A(\hash.CA2.f_dash[0] ),
    .B(\hash.CA2.f_dash[1] ),
    .C(\hash.CA2.f_dash[2] ),
    .Y(_06296_));
 sky130_fd_sc_hd__xnor2_1 _17477_ (.A(\hash.CA2.f_dash[3] ),
    .B(_06296_),
    .Y(_06297_));
 sky130_fd_sc_hd__nor2_1 _17478_ (.A(net343),
    .B(_06297_),
    .Y(_00899_));
 sky130_fd_sc_hd__nor2_4 _17479_ (.A(net344),
    .B(\hash.CA2.f_dash[4] ),
    .Y(_12520_));
 sky130_fd_sc_hd__a21oi_2 _17480_ (.A1(\hash.CA2.f_dash[2] ),
    .A2(_13848_),
    .B1(\hash.CA2.f_dash[3] ),
    .Y(_06298_));
 sky130_fd_sc_hd__xnor2_1 _17481_ (.A(\hash.CA2.f_dash[4] ),
    .B(_06298_),
    .Y(_06299_));
 sky130_fd_sc_hd__nand2_1 _17482_ (.A(_06002_),
    .B(_06299_),
    .Y(_00900_));
 sky130_fd_sc_hd__nor2b_4 _17483_ (.A(net343),
    .B_N(\hash.CA2.f_dash[5] ),
    .Y(_12525_));
 sky130_fd_sc_hd__nand3b_1 _17484_ (.A_N(\hash.CA2.f_dash[3] ),
    .B(_06296_),
    .C(_12520_),
    .Y(_06300_));
 sky130_fd_sc_hd__xor2_1 _17485_ (.A(_12525_),
    .B(_06300_),
    .X(_00901_));
 sky130_fd_sc_hd__nand2_8 _17486_ (.A(_06002_),
    .B(\hash.CA2.f_dash[6] ),
    .Y(_12693_));
 sky130_fd_sc_hd__inv_1 _17487_ (.A(_12693_),
    .Y(_12530_));
 sky130_fd_sc_hd__a21boi_2 _17488_ (.A1(_12520_),
    .A2(_06298_),
    .B1_N(_12525_),
    .Y(_06301_));
 sky130_fd_sc_hd__mux2i_1 _17489_ (.A0(_12693_),
    .A1(\hash.CA2.f_dash[6] ),
    .S(_06301_),
    .Y(_00902_));
 sky130_fd_sc_hd__nand2_8 _17490_ (.A(_06002_),
    .B(\hash.CA2.f_dash[7] ),
    .Y(_12702_));
 sky130_fd_sc_hd__inv_6 _17491_ (.A(_12702_),
    .Y(_12535_));
 sky130_fd_sc_hd__nand3_2 _17492_ (.A(\hash.CA2.f_dash[6] ),
    .B(_12525_),
    .C(_06300_),
    .Y(_06302_));
 sky130_fd_sc_hd__xnor2_1 _17493_ (.A(_12535_),
    .B(_06302_),
    .Y(_00903_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1168 ();
 sky130_fd_sc_hd__nor2_4 _17495_ (.A(net345),
    .B(\hash.CA2.f_dash[8] ),
    .Y(_12540_));
 sky130_fd_sc_hd__and3_4 _17496_ (.A(\hash.CA2.f_dash[6] ),
    .B(_06301_),
    .C(_12535_),
    .X(_06304_));
 sky130_fd_sc_hd__xor2_1 _17497_ (.A(_12540_),
    .B(_06304_),
    .X(_00904_));
 sky130_fd_sc_hd__nand2_8 _17498_ (.A(_06002_),
    .B(\hash.CA2.f_dash[9] ),
    .Y(_12715_));
 sky130_fd_sc_hd__inv_6 _17499_ (.A(_12715_),
    .Y(_12545_));
 sky130_fd_sc_hd__nor2_1 _17500_ (.A(_12702_),
    .B(_06302_),
    .Y(_06305_));
 sky130_fd_sc_hd__o21a_1 _17501_ (.A1(\hash.CA2.f_dash[8] ),
    .A2(_06305_),
    .B1(\hash.CA2.f_dash[9] ),
    .X(_06306_));
 sky130_fd_sc_hd__nor3_1 _17502_ (.A(\hash.CA2.f_dash[8] ),
    .B(\hash.CA2.f_dash[9] ),
    .C(_06305_),
    .Y(_06307_));
 sky130_fd_sc_hd__o21ai_0 _17503_ (.A1(_06306_),
    .A2(_06307_),
    .B1(_06002_),
    .Y(_00905_));
 sky130_fd_sc_hd__nor2_4 _17504_ (.A(net345),
    .B(\hash.CA2.f_dash[10] ),
    .Y(_12550_));
 sky130_fd_sc_hd__o21ai_2 _17505_ (.A1(\hash.CA2.f_dash[8] ),
    .A2(_06304_),
    .B1(_12545_),
    .Y(_06308_));
 sky130_fd_sc_hd__mux2_1 _17506_ (.A0(\hash.CA2.f_dash[10] ),
    .A1(_12550_),
    .S(_06308_),
    .X(_00876_));
 sky130_fd_sc_hd__or2_4 _17507_ (.A(net534),
    .B(\hash.CA2.f_dash[11] ),
    .X(_12733_));
 sky130_fd_sc_hd__inv_1 _17508_ (.A(_12733_),
    .Y(_12555_));
 sky130_fd_sc_hd__or3_1 _17509_ (.A(\hash.CA2.f_dash[10] ),
    .B(\hash.CA2.f_dash[11] ),
    .C(_06306_),
    .X(_06309_));
 sky130_fd_sc_hd__o21ai_0 _17510_ (.A1(\hash.CA2.f_dash[10] ),
    .A2(_06306_),
    .B1(\hash.CA2.f_dash[11] ),
    .Y(_06310_));
 sky130_fd_sc_hd__nand3_1 _17511_ (.A(_06002_),
    .B(_06309_),
    .C(_06310_),
    .Y(_00877_));
 sky130_fd_sc_hd__nand2_4 _17512_ (.A(_06002_),
    .B(\hash.CA2.f_dash[12] ),
    .Y(_06311_));
 sky130_fd_sc_hd__inv_4 _17513_ (.A(_06311_),
    .Y(_12560_));
 sky130_fd_sc_hd__nor3_2 _17514_ (.A(net345),
    .B(\hash.CA2.f_dash[10] ),
    .C(\hash.CA2.f_dash[11] ),
    .Y(_06312_));
 sky130_fd_sc_hd__nand2_2 _17515_ (.A(_06308_),
    .B(_06312_),
    .Y(_06313_));
 sky130_fd_sc_hd__xnor2_1 _17516_ (.A(_06311_),
    .B(_06313_),
    .Y(_00878_));
 sky130_fd_sc_hd__inv_6 _17517_ (.A(\hash.CA2.f_dash[13] ),
    .Y(_06314_));
 sky130_fd_sc_hd__nor2_4 _17518_ (.A(net345),
    .B(_06314_),
    .Y(_12565_));
 sky130_fd_sc_hd__nor3_1 _17519_ (.A(\hash.CA2.f_dash[10] ),
    .B(_12702_),
    .C(_06302_),
    .Y(_06315_));
 sky130_fd_sc_hd__o21ai_2 _17520_ (.A1(\hash.CA2.f_dash[8] ),
    .A2(_06315_),
    .B1(\hash.CA2.f_dash[9] ),
    .Y(_06316_));
 sky130_fd_sc_hd__a21oi_2 _17521_ (.A1(_06312_),
    .A2(_06316_),
    .B1(_06311_),
    .Y(_06317_));
 sky130_fd_sc_hd__mux2_1 _17522_ (.A0(_12565_),
    .A1(_06314_),
    .S(_06317_),
    .X(_00879_));
 sky130_fd_sc_hd__nor2_4 _17523_ (.A(net345),
    .B(\hash.CA2.f_dash[14] ),
    .Y(_12570_));
 sky130_fd_sc_hd__and3_4 _17524_ (.A(\hash.CA2.f_dash[12] ),
    .B(_06313_),
    .C(_12565_),
    .X(_06318_));
 sky130_fd_sc_hd__xor2_1 _17525_ (.A(_12570_),
    .B(_06318_),
    .X(_00880_));
 sky130_fd_sc_hd__nor2_2 _17526_ (.A(net534),
    .B(\hash.CA2.f_dash[15] ),
    .Y(_12575_));
 sky130_fd_sc_hd__a21oi_1 _17527_ (.A1(\hash.CA2.f_dash[13] ),
    .A2(_06317_),
    .B1(\hash.CA2.f_dash[14] ),
    .Y(_06319_));
 sky130_fd_sc_hd__xnor2_1 _17528_ (.A(\hash.CA2.f_dash[15] ),
    .B(_06319_),
    .Y(_06320_));
 sky130_fd_sc_hd__nand2_1 _17529_ (.A(_06002_),
    .B(_06320_),
    .Y(_00881_));
 sky130_fd_sc_hd__nor2b_4 _17530_ (.A(net342),
    .B_N(\hash.CA2.f_dash[16] ),
    .Y(_12580_));
 sky130_fd_sc_hd__nor3_2 _17531_ (.A(net345),
    .B(\hash.CA2.f_dash[14] ),
    .C(\hash.CA2.f_dash[15] ),
    .Y(_06321_));
 sky130_fd_sc_hd__nand2b_1 _17532_ (.A_N(_06318_),
    .B(_06321_),
    .Y(_06322_));
 sky130_fd_sc_hd__xor2_1 _17533_ (.A(_12580_),
    .B(_06322_),
    .X(_00882_));
 sky130_fd_sc_hd__nor2b_4 _17534_ (.A(net342),
    .B_N(\hash.CA2.f_dash[17] ),
    .Y(_12585_));
 sky130_fd_sc_hd__a21boi_2 _17535_ (.A1(\hash.CA2.f_dash[13] ),
    .A2(_06317_),
    .B1_N(_06321_),
    .Y(_06323_));
 sky130_fd_sc_hd__nand2b_1 _17536_ (.A_N(_06323_),
    .B(_12580_),
    .Y(_06324_));
 sky130_fd_sc_hd__xnor2_1 _17537_ (.A(_12585_),
    .B(_06324_),
    .Y(_00883_));
 sky130_fd_sc_hd__nor2b_4 _17538_ (.A(net342),
    .B_N(\hash.CA2.f_dash[18] ),
    .Y(_06325_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1167 ();
 sky130_fd_sc_hd__nand2_2 _17540_ (.A(\hash.CA2.f_dash[17] ),
    .B(_12580_),
    .Y(_06326_));
 sky130_fd_sc_hd__nor2b_4 _17541_ (.A(_06326_),
    .B_N(_06322_),
    .Y(_06327_));
 sky130_fd_sc_hd__xor2_1 _17542_ (.A(_06325_),
    .B(_06327_),
    .X(_00884_));
 sky130_fd_sc_hd__nor2b_4 _17543_ (.A(net342),
    .B_N(\hash.CA2.f_dash[19] ),
    .Y(_12595_));
 sky130_fd_sc_hd__nor2_1 _17544_ (.A(_06323_),
    .B(_06326_),
    .Y(_06328_));
 sky130_fd_sc_hd__nand2_1 _17545_ (.A(\hash.CA2.f_dash[18] ),
    .B(_06328_),
    .Y(_06329_));
 sky130_fd_sc_hd__xnor2_1 _17546_ (.A(_12595_),
    .B(_06329_),
    .Y(_00885_));
 sky130_fd_sc_hd__nand2_4 _17547_ (.A(_06002_),
    .B(\hash.CA2.f_dash[20] ),
    .Y(_12794_));
 sky130_fd_sc_hd__inv_4 _17548_ (.A(_12794_),
    .Y(_12600_));
 sky130_fd_sc_hd__nand3_1 _17549_ (.A(\hash.CA2.f_dash[19] ),
    .B(_06325_),
    .C(_06327_),
    .Y(_06330_));
 sky130_fd_sc_hd__xnor2_1 _17550_ (.A(_12600_),
    .B(_06330_),
    .Y(_00886_));
 sky130_fd_sc_hd__nor2_4 _17551_ (.A(net342),
    .B(\hash.CA2.f_dash[21] ),
    .Y(_12605_));
 sky130_fd_sc_hd__inv_2 _17552_ (.A(_12605_),
    .Y(_12803_));
 sky130_fd_sc_hd__nand3_1 _17553_ (.A(\hash.CA2.f_dash[19] ),
    .B(\hash.CA2.f_dash[20] ),
    .C(_06325_),
    .Y(_06331_));
 sky130_fd_sc_hd__or3_4 _17554_ (.A(_06323_),
    .B(_06326_),
    .C(_06331_),
    .X(_06332_));
 sky130_fd_sc_hd__xnor2_1 _17555_ (.A(_12605_),
    .B(_06332_),
    .Y(_00887_));
 sky130_fd_sc_hd__nor2_4 _17556_ (.A(net534),
    .B(\hash.CA2.f_dash[22] ),
    .Y(_12610_));
 sky130_fd_sc_hd__nand2_1 _17557_ (.A(\hash.CA2.f_dash[19] ),
    .B(_06325_),
    .Y(_06333_));
 sky130_fd_sc_hd__nor3_1 _17558_ (.A(\hash.CA2.f_dash[21] ),
    .B(_12794_),
    .C(_06333_),
    .Y(_06334_));
 sky130_fd_sc_hd__nor2_1 _17559_ (.A(_06321_),
    .B(_06331_),
    .Y(_06335_));
 sky130_fd_sc_hd__a31oi_1 _17560_ (.A1(_06318_),
    .A2(_06321_),
    .A3(_06334_),
    .B1(_06335_),
    .Y(_06336_));
 sky130_fd_sc_hd__o21ai_0 _17561_ (.A1(_06326_),
    .A2(_06336_),
    .B1(_12605_),
    .Y(_06337_));
 sky130_fd_sc_hd__xor2_1 _17562_ (.A(_12610_),
    .B(_06337_),
    .X(_00888_));
 sky130_fd_sc_hd__nor2_2 _17563_ (.A(net534),
    .B(\hash.CA2.f_dash[23] ),
    .Y(_12615_));
 sky130_fd_sc_hd__clkinv_2 _17564_ (.A(_12615_),
    .Y(_12819_));
 sky130_fd_sc_hd__nor2_2 _17565_ (.A(\hash.CA2.f_dash[22] ),
    .B(_12803_),
    .Y(_06338_));
 sky130_fd_sc_hd__nand2_1 _17566_ (.A(_06332_),
    .B(_06338_),
    .Y(_06339_));
 sky130_fd_sc_hd__xnor2_1 _17567_ (.A(_12819_),
    .B(_06339_),
    .Y(_00889_));
 sky130_fd_sc_hd__nor2_2 _17568_ (.A(net534),
    .B(\hash.CA2.f_dash[24] ),
    .Y(_12620_));
 sky130_fd_sc_hd__nand4_1 _17569_ (.A(\hash.CA2.f_dash[19] ),
    .B(\hash.CA2.f_dash[20] ),
    .C(_06325_),
    .D(_06327_),
    .Y(_06340_));
 sky130_fd_sc_hd__nand3b_1 _17570_ (.A_N(\hash.CA2.f_dash[23] ),
    .B(_06338_),
    .C(_06340_),
    .Y(_06341_));
 sky130_fd_sc_hd__xor2_1 _17571_ (.A(\hash.CA2.f_dash[24] ),
    .B(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__nand2_1 _17572_ (.A(_06002_),
    .B(_06342_),
    .Y(_00890_));
 sky130_fd_sc_hd__nor2_4 _17573_ (.A(net342),
    .B(\hash.CA2.f_dash[25] ),
    .Y(_12625_));
 sky130_fd_sc_hd__clkinv_1 _17574_ (.A(_12625_),
    .Y(_12835_));
 sky130_fd_sc_hd__nor2_1 _17575_ (.A(\hash.CA2.f_dash[24] ),
    .B(_12819_),
    .Y(_06343_));
 sky130_fd_sc_hd__nand3_1 _17576_ (.A(_06332_),
    .B(_06338_),
    .C(_06343_),
    .Y(_06344_));
 sky130_fd_sc_hd__xnor2_1 _17577_ (.A(_12835_),
    .B(_06344_),
    .Y(_00891_));
 sky130_fd_sc_hd__nor2b_4 _17578_ (.A(net342),
    .B_N(\hash.CA2.f_dash[26] ),
    .Y(_12630_));
 sky130_fd_sc_hd__nand2_1 _17579_ (.A(_06327_),
    .B(_06334_),
    .Y(_06345_));
 sky130_fd_sc_hd__nand4_1 _17580_ (.A(_06338_),
    .B(_12625_),
    .C(_06343_),
    .D(_06345_),
    .Y(_06346_));
 sky130_fd_sc_hd__xor2_1 _17581_ (.A(_12630_),
    .B(_06346_),
    .X(_00892_));
 sky130_fd_sc_hd__nor2_2 _17582_ (.A(net342),
    .B(\hash.CA2.f_dash[27] ),
    .Y(_12635_));
 sky130_fd_sc_hd__inv_1 _17583_ (.A(_12635_),
    .Y(_12850_));
 sky130_fd_sc_hd__nand4_1 _17584_ (.A(_06332_),
    .B(_06338_),
    .C(_12625_),
    .D(_06343_),
    .Y(_06347_));
 sky130_fd_sc_hd__nand2_1 _17585_ (.A(_12630_),
    .B(_06347_),
    .Y(_06348_));
 sky130_fd_sc_hd__mux2_1 _17586_ (.A0(\hash.CA2.f_dash[27] ),
    .A1(_12635_),
    .S(_06348_),
    .X(_00893_));
 sky130_fd_sc_hd__or2_4 _17587_ (.A(net342),
    .B(\hash.CA2.f_dash[28] ),
    .X(_12858_));
 sky130_fd_sc_hd__inv_1 _17588_ (.A(_12858_),
    .Y(_12640_));
 sky130_fd_sc_hd__a21oi_1 _17589_ (.A1(\hash.CA2.f_dash[26] ),
    .A2(_06346_),
    .B1(\hash.CA2.f_dash[27] ),
    .Y(_06349_));
 sky130_fd_sc_hd__xnor2_1 _17590_ (.A(\hash.CA2.f_dash[28] ),
    .B(_06349_),
    .Y(_06350_));
 sky130_fd_sc_hd__nand2_1 _17591_ (.A(_06002_),
    .B(_06350_),
    .Y(_00894_));
 sky130_fd_sc_hd__nand2_2 _17592_ (.A(_06002_),
    .B(\hash.CA2.f_dash[29] ),
    .Y(_06351_));
 sky130_fd_sc_hd__inv_2 _17593_ (.A(_06351_),
    .Y(_12645_));
 sky130_fd_sc_hd__nor2_1 _17594_ (.A(\hash.CA2.f_dash[27] ),
    .B(_12858_),
    .Y(_06352_));
 sky130_fd_sc_hd__nand2_1 _17595_ (.A(_06348_),
    .B(_06352_),
    .Y(_06353_));
 sky130_fd_sc_hd__xnor2_1 _17596_ (.A(_06351_),
    .B(_06353_),
    .Y(_00895_));
 sky130_fd_sc_hd__nor2_4 _17597_ (.A(net342),
    .B(\hash.CA2.f_dash[30] ),
    .Y(_12650_));
 sky130_fd_sc_hd__inv_1 _17598_ (.A(_12650_),
    .Y(_12872_));
 sky130_fd_sc_hd__and3_1 _17599_ (.A(\hash.CA2.f_dash[26] ),
    .B(\hash.CA2.f_dash[29] ),
    .C(_06352_),
    .X(_06354_));
 sky130_fd_sc_hd__nor2_1 _17600_ (.A(_06351_),
    .B(_06352_),
    .Y(_06355_));
 sky130_fd_sc_hd__a21oi_1 _17601_ (.A1(_06346_),
    .A2(_06354_),
    .B1(_06355_),
    .Y(_06356_));
 sky130_fd_sc_hd__xnor2_1 _17602_ (.A(_12650_),
    .B(_06356_),
    .Y(_00897_));
 sky130_fd_sc_hd__a211oi_1 _17603_ (.A1(_06347_),
    .A2(_06354_),
    .B1(_06355_),
    .C1(\hash.CA2.f_dash[30] ),
    .Y(_06357_));
 sky130_fd_sc_hd__xor2_1 _17604_ (.A(\hash.CA2.f_dash[31] ),
    .B(_06357_),
    .X(_06358_));
 sky130_fd_sc_hd__nand2_1 _17605_ (.A(_06002_),
    .B(_06358_),
    .Y(_00898_));
 sky130_fd_sc_hd__xnor2_1 _17606_ (.A(_13849_),
    .B(_12375_),
    .Y(_00865_));
 sky130_fd_sc_hd__o21ai_2 _17607_ (.A1(\hash.CA2.e_dash[0] ),
    .A2(\hash.CA2.e_dash[1] ),
    .B1(\hash.CA2.e_dash[2] ),
    .Y(_06359_));
 sky130_fd_sc_hd__xnor2_2 _17608_ (.A(\hash.CA2.e_dash[3] ),
    .B(_06359_),
    .Y(_06360_));
 sky130_fd_sc_hd__nor2_1 _17609_ (.A(net340),
    .B(_06360_),
    .Y(_00868_));
 sky130_fd_sc_hd__nor2b_2 _17610_ (.A(_13849_),
    .B_N(\hash.CA2.e_dash[2] ),
    .Y(_06361_));
 sky130_fd_sc_hd__o21a_4 _17611_ (.A1(\hash.CA2.e_dash[3] ),
    .A2(_06361_),
    .B1(\hash.CA2.e_dash[4] ),
    .X(_06362_));
 sky130_fd_sc_hd__nor3_1 _17612_ (.A(\hash.CA2.e_dash[3] ),
    .B(\hash.CA2.e_dash[4] ),
    .C(_06361_),
    .Y(_06363_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1166 ();
 sky130_fd_sc_hd__o21ai_2 _17614_ (.A1(_06362_),
    .A2(_06363_),
    .B1(_06002_),
    .Y(_00869_));
 sky130_fd_sc_hd__o21a_1 _17615_ (.A1(\hash.CA2.e_dash[0] ),
    .A2(\hash.CA2.e_dash[1] ),
    .B1(_12375_),
    .X(_06365_));
 sky130_fd_sc_hd__o21a_4 _17616_ (.A1(\hash.CA2.e_dash[3] ),
    .A2(_06365_),
    .B1(\hash.CA2.e_dash[4] ),
    .X(_06366_));
 sky130_fd_sc_hd__xor2_1 _17617_ (.A(\hash.CA2.e_dash[5] ),
    .B(_06366_),
    .X(_06367_));
 sky130_fd_sc_hd__nor2_1 _17618_ (.A(net343),
    .B(_06367_),
    .Y(_00870_));
 sky130_fd_sc_hd__nor3_1 _17619_ (.A(net343),
    .B(\hash.CA2.e_dash[5] ),
    .C(_06362_),
    .Y(_06368_));
 sky130_fd_sc_hd__xnor2_1 _17620_ (.A(_12394_),
    .B(_06368_),
    .Y(_00871_));
 sky130_fd_sc_hd__o21ai_2 _17621_ (.A1(\hash.CA2.e_dash[5] ),
    .A2(_06366_),
    .B1(\hash.CA2.e_dash[6] ),
    .Y(_06369_));
 sky130_fd_sc_hd__xnor2_1 _17622_ (.A(\hash.CA2.e_dash[7] ),
    .B(_06369_),
    .Y(_06370_));
 sky130_fd_sc_hd__nor2_1 _17623_ (.A(net343),
    .B(_06370_),
    .Y(_00872_));
 sky130_fd_sc_hd__o21ai_2 _17624_ (.A1(\hash.CA2.e_dash[5] ),
    .A2(_06362_),
    .B1(\hash.CA2.e_dash[6] ),
    .Y(_06371_));
 sky130_fd_sc_hd__nand2b_1 _17625_ (.A_N(\hash.CA2.e_dash[7] ),
    .B(_06371_),
    .Y(_06372_));
 sky130_fd_sc_hd__xor2_1 _17626_ (.A(\hash.CA2.e_dash[8] ),
    .B(_06372_),
    .X(_06373_));
 sky130_fd_sc_hd__nand2_1 _17627_ (.A(_06002_),
    .B(_06373_),
    .Y(_00873_));
 sky130_fd_sc_hd__nor3_1 _17628_ (.A(net343),
    .B(\hash.CA2.e_dash[7] ),
    .C(\hash.CA2.e_dash[8] ),
    .Y(_06374_));
 sky130_fd_sc_hd__nand2_1 _17629_ (.A(_06369_),
    .B(_06374_),
    .Y(_06375_));
 sky130_fd_sc_hd__xor2_1 _17630_ (.A(_12407_),
    .B(_06375_),
    .X(_00874_));
 sky130_fd_sc_hd__o21ai_0 _17631_ (.A1(\hash.CA2.e_dash[8] ),
    .A2(_06372_),
    .B1(\hash.CA2.e_dash[9] ),
    .Y(_06376_));
 sky130_fd_sc_hd__xor2_1 _17632_ (.A(\hash.CA2.e_dash[10] ),
    .B(_06376_),
    .X(_06377_));
 sky130_fd_sc_hd__nor2_1 _17633_ (.A(net341),
    .B(_06377_),
    .Y(_00844_));
 sky130_fd_sc_hd__and2_4 _17634_ (.A(\hash.CA2.e_dash[9] ),
    .B(_06375_),
    .X(_06378_));
 sky130_fd_sc_hd__nand2_1 _17635_ (.A(\hash.CA2.e_dash[10] ),
    .B(_06378_),
    .Y(_06379_));
 sky130_fd_sc_hd__xnor2_1 _17636_ (.A(\hash.CA2.e_dash[11] ),
    .B(_06379_),
    .Y(_06380_));
 sky130_fd_sc_hd__nor2_1 _17637_ (.A(net341),
    .B(_06380_),
    .Y(_00845_));
 sky130_fd_sc_hd__nand2_1 _17638_ (.A(\hash.CA2.e_dash[10] ),
    .B(_12407_),
    .Y(_06381_));
 sky130_fd_sc_hd__a21oi_2 _17639_ (.A1(_06371_),
    .A2(_06374_),
    .B1(_06381_),
    .Y(_06382_));
 sky130_fd_sc_hd__or3_1 _17640_ (.A(\hash.CA2.e_dash[11] ),
    .B(\hash.CA2.e_dash[12] ),
    .C(_06382_),
    .X(_06383_));
 sky130_fd_sc_hd__o21ai_0 _17641_ (.A1(\hash.CA2.e_dash[11] ),
    .A2(_06382_),
    .B1(\hash.CA2.e_dash[12] ),
    .Y(_06384_));
 sky130_fd_sc_hd__nand3_1 _17642_ (.A(_06002_),
    .B(_06383_),
    .C(_06384_),
    .Y(_00846_));
 sky130_fd_sc_hd__a211o_1 _17643_ (.A1(_12410_),
    .A2(_06378_),
    .B1(\hash.CA2.e_dash[11] ),
    .C1(\hash.CA2.e_dash[12] ),
    .X(_06385_));
 sky130_fd_sc_hd__or2_0 _17644_ (.A(\hash.CA2.e_dash[13] ),
    .B(_06385_),
    .X(_06386_));
 sky130_fd_sc_hd__nand2_2 _17645_ (.A(\hash.CA2.e_dash[13] ),
    .B(_06385_),
    .Y(_06387_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1165 ();
 sky130_fd_sc_hd__a21o_1 _17647_ (.A1(_06386_),
    .A2(_06387_),
    .B1(net343),
    .X(_00847_));
 sky130_fd_sc_hd__o311a_4 _17648_ (.A1(\hash.CA2.e_dash[11] ),
    .A2(\hash.CA2.e_dash[12] ),
    .A3(_06382_),
    .B1(\hash.CA2.e_dash[13] ),
    .C1(_06002_),
    .X(_06389_));
 sky130_fd_sc_hd__xor2_1 _17649_ (.A(_12428_),
    .B(_06389_),
    .X(_00848_));
 sky130_fd_sc_hd__nand2_1 _17650_ (.A(_12428_),
    .B(_06387_),
    .Y(_06390_));
 sky130_fd_sc_hd__xor2_1 _17651_ (.A(_12433_),
    .B(_06390_),
    .X(_00849_));
 sky130_fd_sc_hd__nor4_1 _17652_ (.A(net343),
    .B(\hash.CA2.e_dash[14] ),
    .C(\hash.CA2.e_dash[15] ),
    .D(_06389_),
    .Y(_06391_));
 sky130_fd_sc_hd__xnor2_1 _17653_ (.A(_12438_),
    .B(_06391_),
    .Y(_00850_));
 sky130_fd_sc_hd__nor4_1 _17654_ (.A(net343),
    .B(\hash.CA2.e_dash[14] ),
    .C(\hash.CA2.e_dash[15] ),
    .D(\hash.CA2.e_dash[16] ),
    .Y(_06392_));
 sky130_fd_sc_hd__nand2_2 _17655_ (.A(_06387_),
    .B(_06392_),
    .Y(_06393_));
 sky130_fd_sc_hd__xor2_1 _17656_ (.A(_12443_),
    .B(_06393_),
    .X(_00851_));
 sky130_fd_sc_hd__or3b_4 _17657_ (.A(\hash.CA2.e_dash[17] ),
    .B(_06389_),
    .C_N(_06392_),
    .X(_06394_));
 sky130_fd_sc_hd__xor2_1 _17658_ (.A(_12446_),
    .B(_06394_),
    .X(_00852_));
 sky130_fd_sc_hd__o31a_1 _17659_ (.A1(net343),
    .A2(\hash.CA2.e_dash[17] ),
    .A3(_06393_),
    .B1(_12446_),
    .X(_06395_));
 sky130_fd_sc_hd__mux2_1 _17660_ (.A0(_12449_),
    .A1(_06294_),
    .S(_06395_),
    .X(_00853_));
 sky130_fd_sc_hd__and3_4 _17661_ (.A(\hash.CA2.e_dash[19] ),
    .B(_12446_),
    .C(_06394_),
    .X(_06396_));
 sky130_fd_sc_hd__xor2_1 _17662_ (.A(_12452_),
    .B(_06396_),
    .X(_00855_));
 sky130_fd_sc_hd__and3_4 _17663_ (.A(\hash.CA2.e_dash[19] ),
    .B(\hash.CA2.e_dash[20] ),
    .C(_06395_),
    .X(_06397_));
 sky130_fd_sc_hd__xor2_1 _17664_ (.A(_12455_),
    .B(_06397_),
    .X(_00856_));
 sky130_fd_sc_hd__nand3_1 _17665_ (.A(\hash.CA2.e_dash[20] ),
    .B(\hash.CA2.e_dash[21] ),
    .C(_06396_),
    .Y(_06398_));
 sky130_fd_sc_hd__xor2_1 _17666_ (.A(\hash.CA2.e_dash[22] ),
    .B(_06398_),
    .X(_06399_));
 sky130_fd_sc_hd__nor2_1 _17667_ (.A(net343),
    .B(_06399_),
    .Y(_00857_));
 sky130_fd_sc_hd__and3_4 _17668_ (.A(\hash.CA2.e_dash[21] ),
    .B(\hash.CA2.e_dash[22] ),
    .C(_12452_),
    .X(_06400_));
 sky130_fd_sc_hd__and3_4 _17669_ (.A(_12449_),
    .B(_06395_),
    .C(_06400_),
    .X(_06401_));
 sky130_fd_sc_hd__xor2_1 _17670_ (.A(_12463_),
    .B(_06401_),
    .X(_00858_));
 sky130_fd_sc_hd__and3_4 _17671_ (.A(_12463_),
    .B(_06396_),
    .C(_06400_),
    .X(_06402_));
 sky130_fd_sc_hd__or3_1 _17672_ (.A(\hash.CA2.e_dash[23] ),
    .B(\hash.CA2.e_dash[24] ),
    .C(_06402_),
    .X(_06403_));
 sky130_fd_sc_hd__o21ai_0 _17673_ (.A1(\hash.CA2.e_dash[23] ),
    .A2(_06402_),
    .B1(\hash.CA2.e_dash[24] ),
    .Y(_06404_));
 sky130_fd_sc_hd__nand3_1 _17674_ (.A(_06002_),
    .B(_06403_),
    .C(_06404_),
    .Y(_00859_));
 sky130_fd_sc_hd__nor3_1 _17675_ (.A(\hash.CA2.e_dash[23] ),
    .B(\hash.CA2.e_dash[24] ),
    .C(_06401_),
    .Y(_06405_));
 sky130_fd_sc_hd__xnor2_1 _17676_ (.A(\hash.CA2.e_dash[25] ),
    .B(_06405_),
    .Y(_06406_));
 sky130_fd_sc_hd__nand2_1 _17677_ (.A(_06002_),
    .B(_06406_),
    .Y(_00860_));
 sky130_fd_sc_hd__nor4_1 _17678_ (.A(\hash.CA2.e_dash[23] ),
    .B(\hash.CA2.e_dash[24] ),
    .C(\hash.CA2.e_dash[25] ),
    .D(_06402_),
    .Y(_06407_));
 sky130_fd_sc_hd__xnor2_1 _17679_ (.A(\hash.CA2.e_dash[26] ),
    .B(_06407_),
    .Y(_06408_));
 sky130_fd_sc_hd__nand2_1 _17680_ (.A(_06002_),
    .B(_06408_),
    .Y(_00861_));
 sky130_fd_sc_hd__nor2_4 _17681_ (.A(\hash.CA2.e_dash[23] ),
    .B(\hash.CA2.e_dash[24] ),
    .Y(_06409_));
 sky130_fd_sc_hd__nor4b_1 _17682_ (.A(\hash.CA2.e_dash[25] ),
    .B(\hash.CA2.e_dash[26] ),
    .C(_06401_),
    .D_N(_06409_),
    .Y(_06410_));
 sky130_fd_sc_hd__xnor2_1 _17683_ (.A(\hash.CA2.e_dash[27] ),
    .B(_06410_),
    .Y(_06411_));
 sky130_fd_sc_hd__nand2_1 _17684_ (.A(_06002_),
    .B(_06411_),
    .Y(_00862_));
 sky130_fd_sc_hd__nand4_1 _17685_ (.A(_12473_),
    .B(_12478_),
    .C(_12483_),
    .D(_06409_),
    .Y(_06412_));
 sky130_fd_sc_hd__nor2_1 _17686_ (.A(_06402_),
    .B(_06412_),
    .Y(_06413_));
 sky130_fd_sc_hd__xnor2_1 _17687_ (.A(_12488_),
    .B(_06413_),
    .Y(_00863_));
 sky130_fd_sc_hd__or2_0 _17688_ (.A(\hash.CA2.e_dash[28] ),
    .B(_06412_),
    .X(_06414_));
 sky130_fd_sc_hd__a41oi_1 _17689_ (.A1(_12455_),
    .A2(_12458_),
    .A3(_06397_),
    .A4(_06409_),
    .B1(_06414_),
    .Y(_06415_));
 sky130_fd_sc_hd__xnor2_1 _17690_ (.A(_12491_),
    .B(_06415_),
    .Y(_00864_));
 sky130_fd_sc_hd__o21ai_1 _17691_ (.A1(_06402_),
    .A2(_06414_),
    .B1(\hash.CA2.e_dash[29] ),
    .Y(_06416_));
 sky130_fd_sc_hd__xor2_1 _17692_ (.A(\hash.CA2.e_dash[30] ),
    .B(_06416_),
    .X(_06417_));
 sky130_fd_sc_hd__nor2_4 _17693_ (.A(net346),
    .B(_06417_),
    .Y(_00866_));
 sky130_fd_sc_hd__nor2b_4 _17694_ (.A(net534),
    .B_N(\hash.CA2.e_dash[31] ),
    .Y(_06418_));
 sky130_fd_sc_hd__nand2_1 _17695_ (.A(\hash.CA2.e_dash[30] ),
    .B(_12491_),
    .Y(_06419_));
 sky130_fd_sc_hd__nor2_1 _17696_ (.A(_06415_),
    .B(_06419_),
    .Y(_06420_));
 sky130_fd_sc_hd__xor2_1 _17697_ (.A(_06418_),
    .B(_06420_),
    .X(_00867_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1164 ();
 sky130_fd_sc_hd__nor2b_1 _17699_ (.A(net344),
    .B_N(\hash.CA2.S1.X[4] ),
    .Y(\hash.CA1.f[4] ));
 sky130_fd_sc_hd__xnor2_1 _17700_ (.A(_13852_),
    .B(\hash.CA1.f[4] ),
    .Y(_00835_));
 sky130_fd_sc_hd__nor2b_1 _17701_ (.A(net343),
    .B_N(\hash.CA2.S1.X[5] ),
    .Y(\hash.CA1.f[5] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1163 ();
 sky130_fd_sc_hd__o21ai_0 _17703_ (.A1(net1121),
    .A2(\hash.CA2.S1.X[3] ),
    .B1(\hash.CA2.S1.X[4] ),
    .Y(_06423_));
 sky130_fd_sc_hd__xor2_1 _17704_ (.A(\hash.CA2.S1.X[5] ),
    .B(_06423_),
    .X(_06424_));
 sky130_fd_sc_hd__nor2_1 _17705_ (.A(net344),
    .B(_06424_),
    .Y(_00836_));
 sky130_fd_sc_hd__nor2b_4 _17706_ (.A(net344),
    .B_N(net1076),
    .Y(\hash.CA1.f[6] ));
 sky130_fd_sc_hd__nor2b_4 _17707_ (.A(_13852_),
    .B_N(\hash.CA2.S1.X[5] ),
    .Y(_06425_));
 sky130_fd_sc_hd__nand2_1 _17708_ (.A(\hash.CA2.S1.X[4] ),
    .B(_06425_),
    .Y(_06426_));
 sky130_fd_sc_hd__xor2_1 _17709_ (.A(net1075),
    .B(_06426_),
    .X(_06427_));
 sky130_fd_sc_hd__nor2_1 _17710_ (.A(net344),
    .B(_06427_),
    .Y(_00837_));
 sky130_fd_sc_hd__clkinv_1 _17711_ (.A(net1084),
    .Y(_06428_));
 sky130_fd_sc_hd__nand2_1 _17712_ (.A(_06002_),
    .B(_06428_),
    .Y(\hash.CA1.f[7] ));
 sky130_fd_sc_hd__o2111ai_2 _17713_ (.A1(net1120),
    .A2(\hash.CA2.S1.X[3] ),
    .B1(\hash.CA2.S1.X[5] ),
    .C1(\hash.CA1.f[4] ),
    .D1(\hash.CA1.f[6] ),
    .Y(_06429_));
 sky130_fd_sc_hd__inv_1 _17714_ (.A(_06429_),
    .Y(_06430_));
 sky130_fd_sc_hd__nand2_1 _17715_ (.A(net1083),
    .B(_06430_),
    .Y(_06431_));
 sky130_fd_sc_hd__o21ai_0 _17716_ (.A1(\hash.CA1.f[7] ),
    .A2(_06430_),
    .B1(_06431_),
    .Y(_00838_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1162 ();
 sky130_fd_sc_hd__clkinvlp_4 _17718_ (.A(net1116),
    .Y(_06433_));
 sky130_fd_sc_hd__nor2_2 _17719_ (.A(net345),
    .B(_06433_),
    .Y(\hash.CA1.f[8] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1161 ();
 sky130_fd_sc_hd__a31oi_4 _17721_ (.A1(net1077),
    .A2(\hash.CA1.f[4] ),
    .A3(_06425_),
    .B1(net1081),
    .Y(_06435_));
 sky130_fd_sc_hd__xnor2_1 _17722_ (.A(_06433_),
    .B(_06435_),
    .Y(_06436_));
 sky130_fd_sc_hd__nand2_1 _17723_ (.A(_06002_),
    .B(_06436_),
    .Y(_00839_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1160 ();
 sky130_fd_sc_hd__nor2b_1 _17725_ (.A(net345),
    .B_N(\hash.CA2.S1.X[9] ),
    .Y(_06438_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1159 ();
 sky130_fd_sc_hd__o21ai_1 _17727_ (.A1(net1081),
    .A2(_06430_),
    .B1(\hash.CA1.f[8] ),
    .Y(_06439_));
 sky130_fd_sc_hd__xnor2_1 _17728_ (.A(_06438_),
    .B(_06439_),
    .Y(_00840_));
 sky130_fd_sc_hd__nor2b_1 _17729_ (.A(net345),
    .B_N(\hash.CA2.S1.X[10] ),
    .Y(\hash.CA1.f[10] ));
 sky130_fd_sc_hd__nand2_1 _17730_ (.A(net1117),
    .B(_06438_),
    .Y(_06440_));
 sky130_fd_sc_hd__nor2_1 _17731_ (.A(_06435_),
    .B(_06440_),
    .Y(_06441_));
 sky130_fd_sc_hd__xor2_1 _17732_ (.A(\hash.CA1.f[10] ),
    .B(_06441_),
    .X(_00841_));
 sky130_fd_sc_hd__nor2_2 _17733_ (.A(net345),
    .B(\hash.CA2.S1.X[11] ),
    .Y(_06442_));
 sky130_fd_sc_hd__clkinvlp_2 _17734_ (.A(_06442_),
    .Y(\hash.CA1.f[11] ));
 sky130_fd_sc_hd__nand2_1 _17735_ (.A(\hash.CA2.S1.X[10] ),
    .B(_06438_),
    .Y(_06443_));
 sky130_fd_sc_hd__nor2_1 _17736_ (.A(_06439_),
    .B(_06443_),
    .Y(_06444_));
 sky130_fd_sc_hd__xnor2_1 _17737_ (.A(\hash.CA1.f[11] ),
    .B(_06444_),
    .Y(_00842_));
 sky130_fd_sc_hd__nor2b_1 _17738_ (.A(net342),
    .B_N(\hash.CA2.S1.X[12] ),
    .Y(\hash.CA1.f[12] ));
 sky130_fd_sc_hd__nand4_1 _17739_ (.A(\hash.CA2.S1.X[8] ),
    .B(\hash.CA2.S1.X[9] ),
    .C(\hash.CA2.S1.X[10] ),
    .D(_06442_),
    .Y(_06445_));
 sky130_fd_sc_hd__nor2_1 _17740_ (.A(_06435_),
    .B(_06445_),
    .Y(_06446_));
 sky130_fd_sc_hd__o21ai_2 _17741_ (.A1(\hash.CA1.f[11] ),
    .A2(_06446_),
    .B1(\hash.CA1.f[12] ),
    .Y(_06447_));
 sky130_fd_sc_hd__o31a_1 _17742_ (.A1(\hash.CA2.S1.X[12] ),
    .A2(\hash.CA1.f[11] ),
    .A3(_06446_),
    .B1(_06447_),
    .X(_00814_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1158 ();
 sky130_fd_sc_hd__or2_0 _17744_ (.A(net345),
    .B(\hash.CA2.S1.X[13] ),
    .X(\hash.CA1.f[13] ));
 sky130_fd_sc_hd__nand2_1 _17745_ (.A(net1082),
    .B(\hash.CA1.f[8] ),
    .Y(_06449_));
 sky130_fd_sc_hd__o32ai_2 _17746_ (.A1(net1082),
    .A2(_06429_),
    .A3(_06445_),
    .B1(_06449_),
    .B2(_06443_),
    .Y(_06450_));
 sky130_fd_sc_hd__o21ai_4 _17747_ (.A1(\hash.CA2.S1.X[11] ),
    .A2(_06450_),
    .B1(\hash.CA1.f[12] ),
    .Y(_06451_));
 sky130_fd_sc_hd__xor2_1 _17748_ (.A(\hash.CA1.f[13] ),
    .B(_06451_),
    .X(_00815_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1157 ();
 sky130_fd_sc_hd__or2_0 _17750_ (.A(net342),
    .B(\hash.CA2.S1.X[14] ),
    .X(\hash.CA1.f[14] ));
 sky130_fd_sc_hd__inv_2 _17751_ (.A(\hash.CA2.S1.X[11] ),
    .Y(_06453_));
 sky130_fd_sc_hd__o21ai_0 _17752_ (.A1(_06435_),
    .A2(_06445_),
    .B1(_06453_),
    .Y(_06454_));
 sky130_fd_sc_hd__a21oi_1 _17753_ (.A1(\hash.CA2.S1.X[12] ),
    .A2(_06454_),
    .B1(\hash.CA2.S1.X[13] ),
    .Y(_06455_));
 sky130_fd_sc_hd__xnor2_1 _17754_ (.A(\hash.CA2.S1.X[14] ),
    .B(_06455_),
    .Y(_06456_));
 sky130_fd_sc_hd__nand2_1 _17755_ (.A(_06002_),
    .B(_06456_),
    .Y(_00816_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1156 ();
 sky130_fd_sc_hd__nand2_2 _17757_ (.A(_06002_),
    .B(\hash.CA2.S1.X[15] ),
    .Y(_06458_));
 sky130_fd_sc_hd__inv_1 _17758_ (.A(_06458_),
    .Y(\hash.CA1.f[15] ));
 sky130_fd_sc_hd__nor2_2 _17759_ (.A(\hash.CA2.S1.X[13] ),
    .B(\hash.CA1.f[14] ),
    .Y(_06459_));
 sky130_fd_sc_hd__nand2_2 _17760_ (.A(_06451_),
    .B(_06459_),
    .Y(_06460_));
 sky130_fd_sc_hd__xnor2_1 _17761_ (.A(_06458_),
    .B(_06460_),
    .Y(_00817_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1155 ();
 sky130_fd_sc_hd__clkinvlp_4 _17763_ (.A(\hash.CA2.S1.X[16] ),
    .Y(_06462_));
 sky130_fd_sc_hd__nand2_2 _17764_ (.A(_06002_),
    .B(_06462_),
    .Y(\hash.CA1.f[16] ));
 sky130_fd_sc_hd__a21oi_2 _17765_ (.A1(_06447_),
    .A2(_06459_),
    .B1(_06458_),
    .Y(_06463_));
 sky130_fd_sc_hd__xnor2_1 _17766_ (.A(\hash.CA1.f[16] ),
    .B(_06463_),
    .Y(_00818_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1154 ();
 sky130_fd_sc_hd__nor2b_1 _17768_ (.A(net342),
    .B_N(\hash.CA2.S1.X[17] ),
    .Y(\hash.CA1.f[17] ));
 sky130_fd_sc_hd__a21o_4 _17769_ (.A1(\hash.CA2.S1.X[15] ),
    .A2(_06460_),
    .B1(\hash.CA1.f[16] ),
    .X(_06465_));
 sky130_fd_sc_hd__xor2_1 _17770_ (.A(\hash.CA1.f[17] ),
    .B(_06465_),
    .X(_00819_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1153 ();
 sky130_fd_sc_hd__or2_0 _17772_ (.A(net342),
    .B(\hash.CA2.S1.X[18] ),
    .X(_06467_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1152 ();
 sky130_fd_sc_hd__o21a_4 _17774_ (.A1(\hash.CA2.S1.X[16] ),
    .A2(_06463_),
    .B1(\hash.CA1.f[17] ),
    .X(_06468_));
 sky130_fd_sc_hd__xnor2_1 _17775_ (.A(_06467_),
    .B(_06468_),
    .Y(_00820_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1151 ();
 sky130_fd_sc_hd__nor2b_1 _17777_ (.A(net342),
    .B_N(\hash.CA2.S1.X[19] ),
    .Y(\hash.CA1.f[19] ));
 sky130_fd_sc_hd__nand2_1 _17778_ (.A(\hash.CA1.f[15] ),
    .B(_06460_),
    .Y(_06470_));
 sky130_fd_sc_hd__nand2_1 _17779_ (.A(_06462_),
    .B(_06470_),
    .Y(_06471_));
 sky130_fd_sc_hd__a21oi_2 _17780_ (.A1(\hash.CA2.S1.X[17] ),
    .A2(_06471_),
    .B1(_06467_),
    .Y(_06472_));
 sky130_fd_sc_hd__xnor2_1 _17781_ (.A(\hash.CA1.f[19] ),
    .B(_06472_),
    .Y(_00821_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1150 ();
 sky130_fd_sc_hd__nor2b_1 _17783_ (.A(net342),
    .B_N(\hash.CA2.S1.X[20] ),
    .Y(\hash.CA1.f[20] ));
 sky130_fd_sc_hd__o21ai_0 _17784_ (.A1(\hash.CA2.S1.X[18] ),
    .A2(_06468_),
    .B1(\hash.CA2.S1.X[19] ),
    .Y(_06474_));
 sky130_fd_sc_hd__xor2_1 _17785_ (.A(\hash.CA2.S1.X[20] ),
    .B(_06474_),
    .X(_06475_));
 sky130_fd_sc_hd__nor2_1 _17786_ (.A(net342),
    .B(_06475_),
    .Y(_00822_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1149 ();
 sky130_fd_sc_hd__nor2b_4 _17788_ (.A(net342),
    .B_N(\hash.CA2.S1.X[21] ),
    .Y(\hash.CA1.f[21] ));
 sky130_fd_sc_hd__nand2_2 _17789_ (.A(\hash.CA2.S1.X[20] ),
    .B(\hash.CA1.f[19] ),
    .Y(_06477_));
 sky130_fd_sc_hd__a21oi_1 _17790_ (.A1(\hash.CA1.f[17] ),
    .A2(_06465_),
    .B1(\hash.CA2.S1.X[18] ),
    .Y(_06478_));
 sky130_fd_sc_hd__nor2_1 _17791_ (.A(_06477_),
    .B(_06478_),
    .Y(_06479_));
 sky130_fd_sc_hd__xor2_1 _17792_ (.A(\hash.CA1.f[21] ),
    .B(_06479_),
    .X(_00823_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1148 ();
 sky130_fd_sc_hd__nor2b_1 _17794_ (.A(net534),
    .B_N(\hash.CA2.S1.X[22] ),
    .Y(\hash.CA1.f[22] ));
 sky130_fd_sc_hd__o2111ai_1 _17795_ (.A1(\hash.CA2.S1.X[18] ),
    .A2(_06468_),
    .B1(\hash.CA1.f[19] ),
    .C1(\hash.CA2.S1.X[20] ),
    .D1(\hash.CA2.S1.X[21] ),
    .Y(_06481_));
 sky130_fd_sc_hd__xor2_1 _17796_ (.A(\hash.CA2.S1.X[22] ),
    .B(_06481_),
    .X(_06482_));
 sky130_fd_sc_hd__nor2_1 _17797_ (.A(net342),
    .B(_06482_),
    .Y(_00825_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1147 ();
 sky130_fd_sc_hd__inv_1 _17799_ (.A(\hash.CA2.S1.X[23] ),
    .Y(_06484_));
 sky130_fd_sc_hd__nor2_1 _17800_ (.A(net342),
    .B(_06484_),
    .Y(\hash.CA1.f[23] ));
 sky130_fd_sc_hd__nand2_2 _17801_ (.A(\hash.CA2.S1.X[22] ),
    .B(\hash.CA1.f[21] ),
    .Y(_06485_));
 sky130_fd_sc_hd__nor3_2 _17802_ (.A(_06472_),
    .B(_06477_),
    .C(_06485_),
    .Y(_06486_));
 sky130_fd_sc_hd__xor2_1 _17803_ (.A(\hash.CA1.f[23] ),
    .B(_06486_),
    .X(_00826_));
 sky130_fd_sc_hd__or2_0 _17804_ (.A(net342),
    .B(\hash.CA2.S1.X[24] ),
    .X(_06487_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1146 ();
 sky130_fd_sc_hd__nor4_1 _17806_ (.A(net342),
    .B(_06484_),
    .C(_06477_),
    .D(_06485_),
    .Y(_06488_));
 sky130_fd_sc_hd__o21ai_1 _17807_ (.A1(_06467_),
    .A2(_06468_),
    .B1(_06488_),
    .Y(_06489_));
 sky130_fd_sc_hd__xor2_1 _17808_ (.A(_06487_),
    .B(_06489_),
    .X(_00827_));
 sky130_fd_sc_hd__clkinvlp_2 _17809_ (.A(net1061),
    .Y(_06490_));
 sky130_fd_sc_hd__nand2_1 _17810_ (.A(_06002_),
    .B(_06490_),
    .Y(\hash.CA1.f[25] ));
 sky130_fd_sc_hd__a21oi_1 _17811_ (.A1(\hash.CA2.S1.X[23] ),
    .A2(_06486_),
    .B1(\hash.CA2.S1.X[24] ),
    .Y(_06491_));
 sky130_fd_sc_hd__xnor2_1 _17812_ (.A(net1060),
    .B(_06491_),
    .Y(_06492_));
 sky130_fd_sc_hd__nand2_1 _17813_ (.A(_06002_),
    .B(_06492_),
    .Y(_00828_));
 sky130_fd_sc_hd__nand2_4 _17814_ (.A(_06002_),
    .B(\hash.CA2.S1.X[26] ),
    .Y(_06493_));
 sky130_fd_sc_hd__inv_1 _17815_ (.A(_06493_),
    .Y(\hash.CA1.f[26] ));
 sky130_fd_sc_hd__nor2_2 _17816_ (.A(net1060),
    .B(_06487_),
    .Y(_06494_));
 sky130_fd_sc_hd__nand2_1 _17817_ (.A(_06489_),
    .B(_06494_),
    .Y(_06495_));
 sky130_fd_sc_hd__xnor2_1 _17818_ (.A(_06493_),
    .B(_06495_),
    .Y(_00829_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1145 ();
 sky130_fd_sc_hd__inv_2 _17820_ (.A(\hash.CA2.S1.X[27] ),
    .Y(_06497_));
 sky130_fd_sc_hd__nand2_1 _17821_ (.A(_06002_),
    .B(_06497_),
    .Y(\hash.CA1.f[27] ));
 sky130_fd_sc_hd__nand2_1 _17822_ (.A(\hash.CA2.S1.X[23] ),
    .B(_06486_),
    .Y(_06498_));
 sky130_fd_sc_hd__a21oi_1 _17823_ (.A1(_06498_),
    .A2(_06494_),
    .B1(_06493_),
    .Y(_06499_));
 sky130_fd_sc_hd__xnor2_1 _17824_ (.A(\hash.CA1.f[27] ),
    .B(_06499_),
    .Y(_00830_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1144 ();
 sky130_fd_sc_hd__inv_4 _17826_ (.A(\hash.CA2.S1.X[28] ),
    .Y(_06501_));
 sky130_fd_sc_hd__nand2_1 _17827_ (.A(_06002_),
    .B(_06501_),
    .Y(\hash.CA1.f[28] ));
 sky130_fd_sc_hd__a21oi_1 _17828_ (.A1(\hash.CA2.S1.X[26] ),
    .A2(_06495_),
    .B1(\hash.CA2.S1.X[27] ),
    .Y(_06502_));
 sky130_fd_sc_hd__xnor2_1 _17829_ (.A(\hash.CA2.S1.X[28] ),
    .B(_06502_),
    .Y(_06503_));
 sky130_fd_sc_hd__nand2_1 _17830_ (.A(_06002_),
    .B(_06503_),
    .Y(_00831_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1143 ();
 sky130_fd_sc_hd__nand2_2 _17832_ (.A(_06002_),
    .B(\hash.CA2.S1.X[29] ),
    .Y(_06505_));
 sky130_fd_sc_hd__inv_1 _17833_ (.A(_06505_),
    .Y(\hash.CA1.f[29] ));
 sky130_fd_sc_hd__nor3_1 _17834_ (.A(_06485_),
    .B(_06487_),
    .C(_06493_),
    .Y(_06506_));
 sky130_fd_sc_hd__nand3_1 _17835_ (.A(\hash.CA2.S1.X[23] ),
    .B(_06479_),
    .C(_06506_),
    .Y(_06507_));
 sky130_fd_sc_hd__nor2_1 _17836_ (.A(\hash.CA2.S1.X[27] ),
    .B(\hash.CA1.f[28] ),
    .Y(_06508_));
 sky130_fd_sc_hd__o211ai_1 _17837_ (.A1(_06493_),
    .A2(_06494_),
    .B1(_06507_),
    .C1(_06508_),
    .Y(_06509_));
 sky130_fd_sc_hd__xnor2_1 _17838_ (.A(_06505_),
    .B(_06509_),
    .Y(_00832_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1142 ();
 sky130_fd_sc_hd__nor2b_1 _17840_ (.A(net534),
    .B_N(\hash.CA2.S1.X[30] ),
    .Y(\hash.CA1.f[30] ));
 sky130_fd_sc_hd__a21oi_1 _17841_ (.A1(_06501_),
    .A2(_06502_),
    .B1(_06505_),
    .Y(_06511_));
 sky130_fd_sc_hd__xor2_1 _17842_ (.A(\hash.CA1.f[30] ),
    .B(_06511_),
    .X(_00833_));
 sky130_fd_sc_hd__or2_0 _17843_ (.A(net534),
    .B(\hash.CA2.S1.X[31] ),
    .X(\hash.CA1.f[31] ));
 sky130_fd_sc_hd__nand3_1 _17844_ (.A(\hash.CA2.S1.X[29] ),
    .B(_06509_),
    .C(\hash.CA1.f[30] ),
    .Y(_06512_));
 sky130_fd_sc_hd__xor2_1 _17845_ (.A(\hash.CA1.f[31] ),
    .B(_06512_),
    .X(_00834_));
 sky130_fd_sc_hd__xor2_2 _17846_ (.A(_12364_),
    .B(_13449_),
    .X(_06513_));
 sky130_fd_sc_hd__nor2_4 _17847_ (.A(net344),
    .B(_06513_),
    .Y(_06514_));
 sky130_fd_sc_hd__inv_4 _17848_ (.A(_06514_),
    .Y(\hash.CA1.S1.X[2] ));
 sky130_fd_sc_hd__xnor2_1 _17849_ (.A(_13855_),
    .B(_06514_),
    .Y(_00803_));
 sky130_fd_sc_hd__nor2_4 _17850_ (.A(net534),
    .B(_12365_),
    .Y(_13854_));
 sky130_fd_sc_hd__clkinvlp_2 _17851_ (.A(_13854_),
    .Y(\hash.CA1.S1.X[1] ));
 sky130_fd_sc_hd__inv_4 _17852_ (.A(_00781_),
    .Y(\hash.CA1.S1.X[0] ));
 sky130_fd_sc_hd__a211oi_2 _17853_ (.A1(_12362_),
    .A2(_13447_),
    .B1(_13446_),
    .C1(_13448_),
    .Y(_06515_));
 sky130_fd_sc_hd__o21ai_2 _17854_ (.A1(_13449_),
    .A2(_13448_),
    .B1(_13451_),
    .Y(_06516_));
 sky130_fd_sc_hd__nor2_4 _17855_ (.A(_06515_),
    .B(_06516_),
    .Y(_06517_));
 sky130_fd_sc_hd__a21o_1 _17856_ (.A1(_12362_),
    .A2(_13447_),
    .B1(_13446_),
    .X(_06518_));
 sky130_fd_sc_hd__a211oi_2 _17857_ (.A1(_13449_),
    .A2(_06518_),
    .B1(_13448_),
    .C1(_13451_),
    .Y(_06519_));
 sky130_fd_sc_hd__o21ai_4 _17858_ (.A1(_06517_),
    .A2(_06519_),
    .B1(_06002_),
    .Y(\hash.CA1.S1.X[3] ));
 sky130_fd_sc_hd__or3_4 _17859_ (.A(_12365_),
    .B(\hash.CA1.S1.X[0] ),
    .C(_06513_),
    .X(_06520_));
 sky130_fd_sc_hd__xnor2_1 _17860_ (.A(\hash.CA1.S1.X[3] ),
    .B(_06520_),
    .Y(_00806_));
 sky130_fd_sc_hd__a21o_1 _17861_ (.A1(_12364_),
    .A2(_13449_),
    .B1(_13448_),
    .X(_06521_));
 sky130_fd_sc_hd__a21oi_4 _17862_ (.A1(_13451_),
    .A2(_06521_),
    .B1(_13450_),
    .Y(_06522_));
 sky130_fd_sc_hd__xnor2_4 _17863_ (.A(_13453_),
    .B(_06522_),
    .Y(_06523_));
 sky130_fd_sc_hd__nor2_4 _17864_ (.A(net344),
    .B(_06523_),
    .Y(_06524_));
 sky130_fd_sc_hd__inv_1 _17865_ (.A(_06524_),
    .Y(\hash.CA1.S1.X[4] ));
 sky130_fd_sc_hd__nand2_1 _17866_ (.A(_13855_),
    .B(_06514_),
    .Y(_06525_));
 sky130_fd_sc_hd__nor2_1 _17867_ (.A(\hash.CA1.S1.X[3] ),
    .B(_06525_),
    .Y(_06526_));
 sky130_fd_sc_hd__xnor2_1 _17868_ (.A(_06524_),
    .B(_06526_),
    .Y(_00807_));
 sky130_fd_sc_hd__o21a_4 _17869_ (.A1(_13453_),
    .A2(_13452_),
    .B1(_13455_),
    .X(_06527_));
 sky130_fd_sc_hd__o31ai_4 _17870_ (.A1(_13450_),
    .A2(_13452_),
    .A3(_06517_),
    .B1(_06527_),
    .Y(_06528_));
 sky130_fd_sc_hd__o21bai_1 _17871_ (.A1(_06515_),
    .A2(_06516_),
    .B1_N(_13450_),
    .Y(_06529_));
 sky130_fd_sc_hd__a211o_4 _17872_ (.A1(_13453_),
    .A2(_06529_),
    .B1(_13452_),
    .C1(_13455_),
    .X(_06530_));
 sky130_fd_sc_hd__a21oi_4 _17873_ (.A1(_06528_),
    .A2(_06530_),
    .B1(net346),
    .Y(_06531_));
 sky130_fd_sc_hd__inv_4 _17874_ (.A(_06531_),
    .Y(\hash.CA1.S1.X[5] ));
 sky130_fd_sc_hd__or3_4 _17875_ (.A(\hash.CA1.S1.X[3] ),
    .B(_06520_),
    .C(_06523_),
    .X(_06532_));
 sky130_fd_sc_hd__xor2_1 _17876_ (.A(_06531_),
    .B(_06532_),
    .X(_00808_));
 sky130_fd_sc_hd__a211oi_2 _17877_ (.A1(_12364_),
    .A2(_13449_),
    .B1(_13448_),
    .C1(_13450_),
    .Y(_06533_));
 sky130_fd_sc_hd__o21ai_2 _17878_ (.A1(_13451_),
    .A2(_13450_),
    .B1(_13453_),
    .Y(_06534_));
 sky130_fd_sc_hd__o21bai_1 _17879_ (.A1(_06533_),
    .A2(_06534_),
    .B1_N(_13452_),
    .Y(_06535_));
 sky130_fd_sc_hd__a21oi_1 _17880_ (.A1(_13455_),
    .A2(_06535_),
    .B1(_13454_),
    .Y(_06536_));
 sky130_fd_sc_hd__xor2_2 _17881_ (.A(_13457_),
    .B(_06536_),
    .X(_06537_));
 sky130_fd_sc_hd__nand2_8 _17882_ (.A(_06002_),
    .B(_06537_),
    .Y(\hash.CA1.S1.X[6] ));
 sky130_fd_sc_hd__nor2_1 _17883_ (.A(\hash.CA1.S1.X[3] ),
    .B(_06523_),
    .Y(_06538_));
 sky130_fd_sc_hd__nand4_1 _17884_ (.A(_13855_),
    .B(_06514_),
    .C(_06531_),
    .D(_06538_),
    .Y(_06539_));
 sky130_fd_sc_hd__xnor2_1 _17885_ (.A(\hash.CA1.S1.X[6] ),
    .B(_06539_),
    .Y(_00809_));
 sky130_fd_sc_hd__nor3_1 _17886_ (.A(_13450_),
    .B(_13452_),
    .C(_13454_),
    .Y(_06540_));
 sky130_fd_sc_hd__o21ai_1 _17887_ (.A1(_06515_),
    .A2(_06516_),
    .B1(_06540_),
    .Y(_06541_));
 sky130_fd_sc_hd__o21a_1 _17888_ (.A1(_13454_),
    .A2(_06527_),
    .B1(_13457_),
    .X(_06542_));
 sky130_fd_sc_hd__a21oi_1 _17889_ (.A1(_06541_),
    .A2(_06542_),
    .B1(_13456_),
    .Y(_06543_));
 sky130_fd_sc_hd__xor2_1 _17890_ (.A(_13459_),
    .B(_06543_),
    .X(_06544_));
 sky130_fd_sc_hd__nor2_4 _17891_ (.A(net346),
    .B(_06544_),
    .Y(\hash.CA1.S1.X[7] ));
 sky130_fd_sc_hd__nor3_1 _17892_ (.A(\hash.CA1.S1.X[5] ),
    .B(_06532_),
    .C(\hash.CA1.S1.X[6] ),
    .Y(_06545_));
 sky130_fd_sc_hd__xnor2_1 _17893_ (.A(\hash.CA1.S1.X[7] ),
    .B(_06545_),
    .Y(_00810_));
 sky130_fd_sc_hd__nor3_1 _17894_ (.A(_13452_),
    .B(_13454_),
    .C(_13456_),
    .Y(_06546_));
 sky130_fd_sc_hd__o21ai_2 _17895_ (.A1(_06533_),
    .A2(_06534_),
    .B1(_06546_),
    .Y(_06547_));
 sky130_fd_sc_hd__o21a_1 _17896_ (.A1(_13455_),
    .A2(_13454_),
    .B1(_13457_),
    .X(_06548_));
 sky130_fd_sc_hd__o21a_1 _17897_ (.A1(_13456_),
    .A2(_06548_),
    .B1(_13459_),
    .X(_06549_));
 sky130_fd_sc_hd__a21oi_2 _17898_ (.A1(_06547_),
    .A2(_06549_),
    .B1(_13458_),
    .Y(_06550_));
 sky130_fd_sc_hd__xnor2_4 _17899_ (.A(net1059),
    .B(_06550_),
    .Y(_06551_));
 sky130_fd_sc_hd__and2_4 _17900_ (.A(_06002_),
    .B(_06551_),
    .X(_06552_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1141 ();
 sky130_fd_sc_hd__o21ai_0 _17902_ (.A1(\hash.CA1.S1.X[6] ),
    .A2(_06539_),
    .B1(\hash.CA1.S1.X[7] ),
    .Y(_06553_));
 sky130_fd_sc_hd__xnor2_1 _17903_ (.A(_06552_),
    .B(_06553_),
    .Y(_00811_));
 sky130_fd_sc_hd__nand4_1 _17904_ (.A(_13459_),
    .B(_13461_),
    .C(_06541_),
    .D(_06542_),
    .Y(_06554_));
 sky130_fd_sc_hd__a21o_1 _17905_ (.A1(_13459_),
    .A2(_13456_),
    .B1(_13458_),
    .X(_06555_));
 sky130_fd_sc_hd__a21oi_1 _17906_ (.A1(_13461_),
    .A2(_06555_),
    .B1(_13460_),
    .Y(_06556_));
 sky130_fd_sc_hd__nand2_4 _17907_ (.A(_06554_),
    .B(_06556_),
    .Y(_06557_));
 sky130_fd_sc_hd__xor2_1 _17908_ (.A(_13463_),
    .B(_06557_),
    .X(_06558_));
 sky130_fd_sc_hd__nor2_4 _17909_ (.A(net346),
    .B(_06558_),
    .Y(_06559_));
 sky130_fd_sc_hd__inv_6 _17910_ (.A(_06559_),
    .Y(\hash.CA1.S1.X[9] ));
 sky130_fd_sc_hd__o311ai_2 _17911_ (.A1(\hash.CA1.S1.X[5] ),
    .A2(_06532_),
    .A3(\hash.CA1.S1.X[6] ),
    .B1(\hash.CA1.S1.X[7] ),
    .C1(_06551_),
    .Y(_06560_));
 sky130_fd_sc_hd__xnor2_1 _17912_ (.A(_06559_),
    .B(_06560_),
    .Y(_00812_));
 sky130_fd_sc_hd__o211ai_1 _17913_ (.A1(\hash.CA1.S1.X[6] ),
    .A2(_06539_),
    .B1(\hash.CA1.S1.X[7] ),
    .C1(_06551_),
    .Y(_06561_));
 sky130_fd_sc_hd__and4_4 _17914_ (.A(_13463_),
    .B(_13461_),
    .C(_06547_),
    .D(_06549_),
    .X(_06562_));
 sky130_fd_sc_hd__a21o_1 _17915_ (.A1(_13461_),
    .A2(_13458_),
    .B1(_13460_),
    .X(_06563_));
 sky130_fd_sc_hd__a21oi_2 _17916_ (.A1(_13463_),
    .A2(_06563_),
    .B1(_13462_),
    .Y(_06564_));
 sky130_fd_sc_hd__clkinv_2 _17917_ (.A(_06564_),
    .Y(_06565_));
 sky130_fd_sc_hd__nor2_2 _17918_ (.A(_06562_),
    .B(_06565_),
    .Y(_06566_));
 sky130_fd_sc_hd__xnor2_2 _17919_ (.A(_13465_),
    .B(_06566_),
    .Y(_06567_));
 sky130_fd_sc_hd__nand2_8 _17920_ (.A(_06002_),
    .B(_06567_),
    .Y(_06568_));
 sky130_fd_sc_hd__a21oi_2 _17921_ (.A1(_06559_),
    .A2(_06561_),
    .B1(_06568_),
    .Y(_06569_));
 sky130_fd_sc_hd__and3_1 _17922_ (.A(_06559_),
    .B(_06568_),
    .C(_06561_),
    .X(_06570_));
 sky130_fd_sc_hd__nor2_1 _17923_ (.A(_06569_),
    .B(_06570_),
    .Y(_00782_));
 sky130_fd_sc_hd__nor2_1 _17924_ (.A(net346),
    .B(_13467_),
    .Y(_06571_));
 sky130_fd_sc_hd__nor2b_1 _17925_ (.A(net346),
    .B_N(_13467_),
    .Y(_06572_));
 sky130_fd_sc_hd__a21o_1 _17926_ (.A1(_13463_),
    .A2(_06557_),
    .B1(_13462_),
    .X(_06573_));
 sky130_fd_sc_hd__a21oi_1 _17927_ (.A1(_13465_),
    .A2(_06573_),
    .B1(_13464_),
    .Y(_06574_));
 sky130_fd_sc_hd__mux2_8 _17928_ (.A0(_06571_),
    .A1(_06572_),
    .S(_06574_),
    .X(_06575_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1140 ();
 sky130_fd_sc_hd__a21oi_4 _17930_ (.A1(_06559_),
    .A2(_06560_),
    .B1(_06568_),
    .Y(_06576_));
 sky130_fd_sc_hd__xor2_1 _17931_ (.A(_06575_),
    .B(_06576_),
    .X(_00783_));
 sky130_fd_sc_hd__a21o_4 _17932_ (.A1(_13467_),
    .A2(_13464_),
    .B1(_13466_),
    .X(_06577_));
 sky130_fd_sc_hd__o211a_1 _17933_ (.A1(_06562_),
    .A2(_06565_),
    .B1(_13465_),
    .C1(_13467_),
    .X(_06578_));
 sky130_fd_sc_hd__nor2_1 _17934_ (.A(_06577_),
    .B(_06578_),
    .Y(_06579_));
 sky130_fd_sc_hd__xnor2_1 _17935_ (.A(_13469_),
    .B(_06579_),
    .Y(_06580_));
 sky130_fd_sc_hd__nor2_4 _17936_ (.A(net346),
    .B(_06580_),
    .Y(_06581_));
 sky130_fd_sc_hd__inv_2 _17937_ (.A(_06581_),
    .Y(\hash.CA1.S1.X[12] ));
 sky130_fd_sc_hd__nand2_1 _17938_ (.A(_06569_),
    .B(_06575_),
    .Y(_06582_));
 sky130_fd_sc_hd__xnor2_1 _17939_ (.A(_06581_),
    .B(_06582_),
    .Y(_00784_));
 sky130_fd_sc_hd__nor2_1 _17940_ (.A(net346),
    .B(_13471_),
    .Y(_06583_));
 sky130_fd_sc_hd__nor2b_2 _17941_ (.A(net346),
    .B_N(_13471_),
    .Y(_06584_));
 sky130_fd_sc_hd__a21oi_1 _17942_ (.A1(_13463_),
    .A2(_06557_),
    .B1(_13462_),
    .Y(_06585_));
 sky130_fd_sc_hd__nand3_2 _17943_ (.A(_13469_),
    .B(_13465_),
    .C(_13467_),
    .Y(_06586_));
 sky130_fd_sc_hd__a21oi_4 _17944_ (.A1(_06577_),
    .A2(_13469_),
    .B1(_13468_),
    .Y(_06587_));
 sky130_fd_sc_hd__o21a_4 _17945_ (.A1(_06585_),
    .A2(_06586_),
    .B1(_06587_),
    .X(_06588_));
 sky130_fd_sc_hd__mux2i_4 _17946_ (.A0(_06583_),
    .A1(_06584_),
    .S(_06588_),
    .Y(_06589_));
 sky130_fd_sc_hd__inv_8 _17947_ (.A(_06589_),
    .Y(\hash.CA1.S1.X[13] ));
 sky130_fd_sc_hd__nand2_1 _17948_ (.A(_06575_),
    .B(_06576_),
    .Y(_06590_));
 sky130_fd_sc_hd__nand2_1 _17949_ (.A(_06581_),
    .B(_06590_),
    .Y(_06591_));
 sky130_fd_sc_hd__xnor2_1 _17950_ (.A(_06589_),
    .B(_06591_),
    .Y(_00785_));
 sky130_fd_sc_hd__o211a_1 _17951_ (.A1(_06577_),
    .A2(_06578_),
    .B1(_13469_),
    .C1(_13471_),
    .X(_06592_));
 sky130_fd_sc_hd__a21oi_1 _17952_ (.A1(_13471_),
    .A2(_13468_),
    .B1(_13470_),
    .Y(_06593_));
 sky130_fd_sc_hd__inv_1 _17953_ (.A(_06593_),
    .Y(_06594_));
 sky130_fd_sc_hd__o21ai_2 _17954_ (.A1(_06592_),
    .A2(_06594_),
    .B1(_13473_),
    .Y(_06595_));
 sky130_fd_sc_hd__or3_4 _17955_ (.A(_13473_),
    .B(_06592_),
    .C(_06594_),
    .X(_06596_));
 sky130_fd_sc_hd__a21oi_4 _17956_ (.A1(_06595_),
    .A2(_06596_),
    .B1(net346),
    .Y(_06597_));
 sky130_fd_sc_hd__inv_4 _17957_ (.A(_06597_),
    .Y(\hash.CA1.S1.X[14] ));
 sky130_fd_sc_hd__a21boi_2 _17958_ (.A1(_06569_),
    .A2(_06575_),
    .B1_N(_06581_),
    .Y(_06598_));
 sky130_fd_sc_hd__nand2_1 _17959_ (.A(\hash.CA1.S1.X[13] ),
    .B(\hash.CA1.S1.X[14] ),
    .Y(_06599_));
 sky130_fd_sc_hd__o21ai_4 _17960_ (.A1(_06598_),
    .A2(_06589_),
    .B1(_06597_),
    .Y(_06600_));
 sky130_fd_sc_hd__o21ai_0 _17961_ (.A1(_06598_),
    .A2(_06599_),
    .B1(_06600_),
    .Y(_00786_));
 sky130_fd_sc_hd__nand2_2 _17962_ (.A(_13473_),
    .B(_13471_),
    .Y(_06601_));
 sky130_fd_sc_hd__a21oi_2 _17963_ (.A1(_13470_),
    .A2(_13473_),
    .B1(_13472_),
    .Y(_06602_));
 sky130_fd_sc_hd__o21ai_2 _17964_ (.A1(_06587_),
    .A2(_06601_),
    .B1(_06602_),
    .Y(_06603_));
 sky130_fd_sc_hd__o21a_1 _17965_ (.A1(_06587_),
    .A2(_06601_),
    .B1(_06602_),
    .X(_06604_));
 sky130_fd_sc_hd__nor2_1 _17966_ (.A(_06586_),
    .B(_06601_),
    .Y(_06605_));
 sky130_fd_sc_hd__o21ai_0 _17967_ (.A1(_13463_),
    .A2(_13462_),
    .B1(_06605_),
    .Y(_06606_));
 sky130_fd_sc_hd__nand2_1 _17968_ (.A(_06604_),
    .B(_06606_),
    .Y(_06607_));
 sky130_fd_sc_hd__o31a_1 _17969_ (.A1(_13462_),
    .A2(_06557_),
    .A3(_06603_),
    .B1(_06607_),
    .X(_06608_));
 sky130_fd_sc_hd__xnor2_1 _17970_ (.A(_13475_),
    .B(_06608_),
    .Y(_06609_));
 sky130_fd_sc_hd__nor2_4 _17971_ (.A(net346),
    .B(_06609_),
    .Y(_06610_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1139 ();
 sky130_fd_sc_hd__o21a_1 _17973_ (.A1(_06581_),
    .A2(_06589_),
    .B1(_06597_),
    .X(_06611_));
 sky130_fd_sc_hd__nand3_1 _17974_ (.A(_06575_),
    .B(_06576_),
    .C(\hash.CA1.S1.X[13] ),
    .Y(_06612_));
 sky130_fd_sc_hd__nand2_1 _17975_ (.A(_06611_),
    .B(_06612_),
    .Y(_06613_));
 sky130_fd_sc_hd__xor2_1 _17976_ (.A(_06610_),
    .B(_06613_),
    .X(_00787_));
 sky130_fd_sc_hd__nor2_1 _17977_ (.A(_13474_),
    .B(_06605_),
    .Y(_06614_));
 sky130_fd_sc_hd__nor2_1 _17978_ (.A(_13475_),
    .B(_13474_),
    .Y(_06615_));
 sky130_fd_sc_hd__a21oi_1 _17979_ (.A1(_06604_),
    .A2(_06614_),
    .B1(_06615_),
    .Y(_06616_));
 sky130_fd_sc_hd__or4_4 _17980_ (.A(_13474_),
    .B(_06562_),
    .C(_06565_),
    .D(_06603_),
    .X(_06617_));
 sky130_fd_sc_hd__and2_4 _17981_ (.A(_06616_),
    .B(_06617_),
    .X(_06618_));
 sky130_fd_sc_hd__xnor2_1 _17982_ (.A(_13477_),
    .B(_06618_),
    .Y(_06619_));
 sky130_fd_sc_hd__nor2_4 _17983_ (.A(net346),
    .B(_06619_),
    .Y(\hash.CA1.S1.X[16] ));
 sky130_fd_sc_hd__nand2_1 _17984_ (.A(_06600_),
    .B(_06610_),
    .Y(_06620_));
 sky130_fd_sc_hd__xnor2_1 _17985_ (.A(\hash.CA1.S1.X[16] ),
    .B(_06620_),
    .Y(_00788_));
 sky130_fd_sc_hd__a21o_1 _17986_ (.A1(_13477_),
    .A2(_13474_),
    .B1(_13476_),
    .X(_06621_));
 sky130_fd_sc_hd__a31oi_1 _17987_ (.A1(_13475_),
    .A2(_13481_),
    .A3(_06608_),
    .B1(_06621_),
    .Y(_06622_));
 sky130_fd_sc_hd__xnor2_1 _17988_ (.A(_13479_),
    .B(_06622_),
    .Y(_06623_));
 sky130_fd_sc_hd__nor2_4 _17989_ (.A(\hash.reset ),
    .B(_06623_),
    .Y(_06624_));
 sky130_fd_sc_hd__inv_1 _17990_ (.A(_06624_),
    .Y(\hash.CA1.S1.X[17] ));
 sky130_fd_sc_hd__nand2_1 _17991_ (.A(_06610_),
    .B(\hash.CA1.S1.X[16] ),
    .Y(_06625_));
 sky130_fd_sc_hd__a21o_4 _17992_ (.A1(_06611_),
    .A2(_06612_),
    .B1(_06625_),
    .X(_06626_));
 sky130_fd_sc_hd__xnor2_1 _17993_ (.A(_06624_),
    .B(_06626_),
    .Y(_00789_));
 sky130_fd_sc_hd__a211oi_4 _17994_ (.A1(_06617_),
    .A2(_06616_),
    .B1(_13476_),
    .C1(_13478_),
    .Y(_06627_));
 sky130_fd_sc_hd__o21a_1 _17995_ (.A1(_13481_),
    .A2(_13476_),
    .B1(_13479_),
    .X(_06628_));
 sky130_fd_sc_hd__o21ai_1 _17996_ (.A1(_13478_),
    .A2(_06628_),
    .B1(_13483_),
    .Y(_06629_));
 sky130_fd_sc_hd__or2_4 _17997_ (.A(_06627_),
    .B(_06629_),
    .X(_06630_));
 sky130_fd_sc_hd__o21ai_0 _17998_ (.A1(_13476_),
    .A2(_06618_),
    .B1(_06628_),
    .Y(_06631_));
 sky130_fd_sc_hd__nor2_1 _17999_ (.A(_13483_),
    .B(_13478_),
    .Y(_06632_));
 sky130_fd_sc_hd__nand2_2 _18000_ (.A(_06631_),
    .B(_06632_),
    .Y(_06633_));
 sky130_fd_sc_hd__a21oi_4 _18001_ (.A1(_06630_),
    .A2(_06633_),
    .B1(net346),
    .Y(_06634_));
 sky130_fd_sc_hd__inv_1 _18002_ (.A(_06634_),
    .Y(\hash.CA1.S1.X[18] ));
 sky130_fd_sc_hd__a31oi_1 _18003_ (.A1(_06600_),
    .A2(_06610_),
    .A3(\hash.CA1.S1.X[16] ),
    .B1(\hash.CA1.S1.X[17] ),
    .Y(_06635_));
 sky130_fd_sc_hd__xnor2_1 _18004_ (.A(_06634_),
    .B(_06635_),
    .Y(_00790_));
 sky130_fd_sc_hd__a21o_1 _18005_ (.A1(_13479_),
    .A2(_06621_),
    .B1(_13478_),
    .X(_06636_));
 sky130_fd_sc_hd__a21oi_2 _18006_ (.A1(_13483_),
    .A2(_06636_),
    .B1(_13482_),
    .Y(_06637_));
 sky130_fd_sc_hd__and4_4 _18007_ (.A(_13475_),
    .B(_13479_),
    .C(_13481_),
    .D(_13483_),
    .X(_06638_));
 sky130_fd_sc_hd__o311ai_2 _18008_ (.A1(_13462_),
    .A2(_06557_),
    .A3(_06603_),
    .B1(_06607_),
    .C1(_06638_),
    .Y(_06639_));
 sky130_fd_sc_hd__and2_4 _18009_ (.A(_06637_),
    .B(_06639_),
    .X(_06640_));
 sky130_fd_sc_hd__xnor2_1 _18010_ (.A(_13485_),
    .B(_06640_),
    .Y(_06641_));
 sky130_fd_sc_hd__nor2_4 _18011_ (.A(net346),
    .B(_06641_),
    .Y(_06642_));
 sky130_fd_sc_hd__inv_1 _18012_ (.A(_06642_),
    .Y(\hash.CA1.S1.X[19] ));
 sky130_fd_sc_hd__nand3_1 _18013_ (.A(_06624_),
    .B(_06626_),
    .C(_06634_),
    .Y(_06643_));
 sky130_fd_sc_hd__xnor2_1 _18014_ (.A(\hash.CA1.S1.X[19] ),
    .B(_06643_),
    .Y(_00791_));
 sky130_fd_sc_hd__nor2_1 _18015_ (.A(_13482_),
    .B(_13484_),
    .Y(_06644_));
 sky130_fd_sc_hd__or2_0 _18016_ (.A(_13485_),
    .B(_13484_),
    .X(_06645_));
 sky130_fd_sc_hd__a21boi_2 _18017_ (.A1(_06630_),
    .A2(_06644_),
    .B1_N(_06645_),
    .Y(_06646_));
 sky130_fd_sc_hd__xnor2_2 _18018_ (.A(_13487_),
    .B(_06646_),
    .Y(_06647_));
 sky130_fd_sc_hd__nor2_4 _18019_ (.A(net534),
    .B(_06647_),
    .Y(\hash.CA1.S1.X[20] ));
 sky130_fd_sc_hd__nand3_4 _18020_ (.A(_06624_),
    .B(_06634_),
    .C(_06642_),
    .Y(_06648_));
 sky130_fd_sc_hd__a31oi_4 _18021_ (.A1(_06600_),
    .A2(_06610_),
    .A3(\hash.CA1.S1.X[16] ),
    .B1(_06648_),
    .Y(_06649_));
 sky130_fd_sc_hd__xnor2_1 _18022_ (.A(\hash.CA1.S1.X[20] ),
    .B(_06649_),
    .Y(_00793_));
 sky130_fd_sc_hd__nand2_2 _18023_ (.A(_13485_),
    .B(_13491_),
    .Y(_06650_));
 sky130_fd_sc_hd__a21oi_2 _18024_ (.A1(_13487_),
    .A2(_13484_),
    .B1(_13486_),
    .Y(_06651_));
 sky130_fd_sc_hd__o21ai_4 _18025_ (.A1(_06640_),
    .A2(_06650_),
    .B1(_06651_),
    .Y(_06652_));
 sky130_fd_sc_hd__xnor2_4 _18026_ (.A(_13489_),
    .B(_06652_),
    .Y(_06653_));
 sky130_fd_sc_hd__nor2_4 _18027_ (.A(net534),
    .B(_06653_),
    .Y(\hash.CA1.S1.X[21] ));
 sky130_fd_sc_hd__nor2b_4 _18028_ (.A(_06648_),
    .B_N(_06626_),
    .Y(_06654_));
 sky130_fd_sc_hd__nand2b_1 _18029_ (.A_N(_06654_),
    .B(\hash.CA1.S1.X[20] ),
    .Y(_06655_));
 sky130_fd_sc_hd__xnor2_1 _18030_ (.A(\hash.CA1.S1.X[21] ),
    .B(_06655_),
    .Y(_00794_));
 sky130_fd_sc_hd__a21o_1 _18031_ (.A1(_13489_),
    .A2(_13486_),
    .B1(_13488_),
    .X(_06656_));
 sky130_fd_sc_hd__nor3_2 _18032_ (.A(_13482_),
    .B(_06656_),
    .C(_13484_),
    .Y(_06657_));
 sky130_fd_sc_hd__a31oi_2 _18033_ (.A1(_13491_),
    .A2(_13495_),
    .A3(_06645_),
    .B1(_06656_),
    .Y(_06658_));
 sky130_fd_sc_hd__a21oi_1 _18034_ (.A1(_06630_),
    .A2(_06657_),
    .B1(_06658_),
    .Y(_06659_));
 sky130_fd_sc_hd__xnor2_1 _18035_ (.A(_13493_),
    .B(_06659_),
    .Y(_06660_));
 sky130_fd_sc_hd__nor2_4 _18036_ (.A(net346),
    .B(_06660_),
    .Y(\hash.CA1.S1.X[22] ));
 sky130_fd_sc_hd__nor4_1 _18037_ (.A(net534),
    .B(_06647_),
    .C(_06649_),
    .D(_06653_),
    .Y(_06661_));
 sky130_fd_sc_hd__xor2_2 _18038_ (.A(\hash.CA1.S1.X[22] ),
    .B(_06661_),
    .X(_00795_));
 sky130_fd_sc_hd__a21o_4 _18039_ (.A1(_13493_),
    .A2(_13488_),
    .B1(_13492_),
    .X(_06662_));
 sky130_fd_sc_hd__a31oi_4 _18040_ (.A1(_13495_),
    .A2(_13499_),
    .A3(_06652_),
    .B1(_06662_),
    .Y(_06663_));
 sky130_fd_sc_hd__xnor2_4 _18041_ (.A(_13497_),
    .B(_06663_),
    .Y(_06664_));
 sky130_fd_sc_hd__nand2_8 _18042_ (.A(_06002_),
    .B(_06664_),
    .Y(_06665_));
 sky130_fd_sc_hd__inv_6 _18043_ (.A(_06665_),
    .Y(\hash.CA1.S1.X[23] ));
 sky130_fd_sc_hd__nand3_4 _18044_ (.A(\hash.CA1.S1.X[20] ),
    .B(\hash.CA1.S1.X[21] ),
    .C(\hash.CA1.S1.X[22] ),
    .Y(_06666_));
 sky130_fd_sc_hd__nor2_1 _18045_ (.A(_06654_),
    .B(_06666_),
    .Y(_06667_));
 sky130_fd_sc_hd__xnor2_1 _18046_ (.A(_06665_),
    .B(_06667_),
    .Y(_00796_));
 sky130_fd_sc_hd__o21ai_2 _18047_ (.A1(_06629_),
    .A2(_06627_),
    .B1(_06657_),
    .Y(_06668_));
 sky130_fd_sc_hd__nand2_1 _18048_ (.A(_13499_),
    .B(_13503_),
    .Y(_06669_));
 sky130_fd_sc_hd__nor2_2 _18049_ (.A(_06658_),
    .B(_06669_),
    .Y(_06670_));
 sky130_fd_sc_hd__a221oi_4 _18050_ (.A1(_13497_),
    .A2(_13492_),
    .B1(_06668_),
    .B2(_06670_),
    .C1(_13496_),
    .Y(_06671_));
 sky130_fd_sc_hd__xnor2_1 _18051_ (.A(_13501_),
    .B(_06671_),
    .Y(_06672_));
 sky130_fd_sc_hd__nor2_4 _18052_ (.A(net534),
    .B(_06672_),
    .Y(_06673_));
 sky130_fd_sc_hd__inv_1 _18053_ (.A(_06673_),
    .Y(\hash.CA1.S1.X[24] ));
 sky130_fd_sc_hd__o31ai_2 _18054_ (.A1(_06649_),
    .A2(_06665_),
    .A3(_06666_),
    .B1(_06673_),
    .Y(_06674_));
 sky130_fd_sc_hd__or4_1 _18055_ (.A(_06649_),
    .B(_06665_),
    .C(_06666_),
    .D(_06673_),
    .X(_06675_));
 sky130_fd_sc_hd__nand2_1 _18056_ (.A(_06674_),
    .B(_06675_),
    .Y(_00797_));
 sky130_fd_sc_hd__nand3_1 _18057_ (.A(_13495_),
    .B(_13499_),
    .C(_13503_),
    .Y(_06676_));
 sky130_fd_sc_hd__a211oi_2 _18058_ (.A1(_06639_),
    .A2(_06637_),
    .B1(_06650_),
    .C1(_06676_),
    .Y(_06677_));
 sky130_fd_sc_hd__nand2_2 _18059_ (.A(_13503_),
    .B(_06662_),
    .Y(_06678_));
 sky130_fd_sc_hd__o21ai_2 _18060_ (.A1(_06651_),
    .A2(_06676_),
    .B1(_06678_),
    .Y(_06679_));
 sky130_fd_sc_hd__or3_4 _18061_ (.A(_06679_),
    .B(_06677_),
    .C(_13496_),
    .X(_06680_));
 sky130_fd_sc_hd__a21oi_4 _18062_ (.A1(_13501_),
    .A2(_06680_),
    .B1(_13500_),
    .Y(_06681_));
 sky130_fd_sc_hd__xor2_2 _18063_ (.A(_13505_),
    .B(_06681_),
    .X(_06682_));
 sky130_fd_sc_hd__nor2_4 _18064_ (.A(net344),
    .B(_06682_),
    .Y(_06683_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1138 ();
 sky130_fd_sc_hd__o31ai_4 _18066_ (.A1(_06654_),
    .A2(_06665_),
    .A3(_06666_),
    .B1(_06673_),
    .Y(_06684_));
 sky130_fd_sc_hd__xor2_1 _18067_ (.A(net1054),
    .B(_06684_),
    .X(_00798_));
 sky130_fd_sc_hd__nand2_1 _18068_ (.A(_13501_),
    .B(_13509_),
    .Y(_06685_));
 sky130_fd_sc_hd__a21oi_1 _18069_ (.A1(_13505_),
    .A2(_13500_),
    .B1(_13504_),
    .Y(_06686_));
 sky130_fd_sc_hd__o21ai_1 _18070_ (.A1(_06671_),
    .A2(_06685_),
    .B1(_06686_),
    .Y(_06687_));
 sky130_fd_sc_hd__xnor2_1 _18071_ (.A(_06687_),
    .B(_13507_),
    .Y(_06688_));
 sky130_fd_sc_hd__nor2_4 _18072_ (.A(_06688_),
    .B(net345),
    .Y(_06689_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1137 ();
 sky130_fd_sc_hd__nand2_1 _18074_ (.A(_06674_),
    .B(net1054),
    .Y(_06690_));
 sky130_fd_sc_hd__xnor2_2 _18075_ (.A(net1057),
    .B(_06690_),
    .Y(_00799_));
 sky130_fd_sc_hd__a21o_4 _18076_ (.A1(_13507_),
    .A2(_13504_),
    .B1(_13506_),
    .X(_06691_));
 sky130_fd_sc_hd__or3_1 _18077_ (.A(_13496_),
    .B(_13500_),
    .C(_06691_),
    .X(_06692_));
 sky130_fd_sc_hd__or3_4 _18078_ (.A(_06677_),
    .B(_06679_),
    .C(_06692_),
    .X(_06693_));
 sky130_fd_sc_hd__a21oi_1 _18079_ (.A1(_13509_),
    .A2(_13513_),
    .B1(_06691_),
    .Y(_06694_));
 sky130_fd_sc_hd__nor3_1 _18080_ (.A(_13501_),
    .B(_13500_),
    .C(_06691_),
    .Y(_06695_));
 sky130_fd_sc_hd__nor2_1 _18081_ (.A(_06694_),
    .B(_06695_),
    .Y(_06696_));
 sky130_fd_sc_hd__nand2_1 _18082_ (.A(_06693_),
    .B(_06696_),
    .Y(_06697_));
 sky130_fd_sc_hd__xor2_1 _18083_ (.A(_13511_),
    .B(_06697_),
    .X(_06698_));
 sky130_fd_sc_hd__nor2_4 _18084_ (.A(_06698_),
    .B(net534),
    .Y(_06699_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1136 ();
 sky130_fd_sc_hd__nand3_2 _18086_ (.A(net1054),
    .B(_06684_),
    .C(net1056),
    .Y(_06700_));
 sky130_fd_sc_hd__xnor2_2 _18087_ (.A(net1124),
    .B(_06700_),
    .Y(_00800_));
 sky130_fd_sc_hd__nor2b_1 _18088_ (.A(_06686_),
    .B_N(_13507_),
    .Y(_06701_));
 sky130_fd_sc_hd__nand3_1 _18089_ (.A(_13507_),
    .B(_13501_),
    .C(_13509_),
    .Y(_06702_));
 sky130_fd_sc_hd__nor2_2 _18090_ (.A(_06702_),
    .B(_06671_),
    .Y(_06703_));
 sky130_fd_sc_hd__o31a_1 _18091_ (.A1(_13506_),
    .A2(_06701_),
    .A3(_06703_),
    .B1(_13511_),
    .X(_06704_));
 sky130_fd_sc_hd__o21ai_4 _18092_ (.A1(_13510_),
    .A2(_06704_),
    .B1(_13515_),
    .Y(_06705_));
 sky130_fd_sc_hd__or3_1 _18093_ (.A(net534),
    .B(_13515_),
    .C(_13510_),
    .X(_06706_));
 sky130_fd_sc_hd__o22a_4 _18094_ (.A1(net345),
    .A2(_06705_),
    .B1(_06706_),
    .B2(_06704_),
    .X(_06707_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1135 ();
 sky130_fd_sc_hd__nand4_1 _18096_ (.A(_06674_),
    .B(net1054),
    .C(net1057),
    .D(net1124),
    .Y(_06708_));
 sky130_fd_sc_hd__xor2_1 _18097_ (.A(net1097),
    .B(_06708_),
    .X(_00801_));
 sky130_fd_sc_hd__a31o_4 _18098_ (.A1(_06693_),
    .A2(_13511_),
    .A3(_06696_),
    .B1(_13510_),
    .X(_06709_));
 sky130_fd_sc_hd__a21oi_4 _18099_ (.A1(_13515_),
    .A2(_06709_),
    .B1(_13514_),
    .Y(_06710_));
 sky130_fd_sc_hd__xnor2_4 _18100_ (.A(net1123),
    .B(_13517_),
    .Y(_06711_));
 sky130_fd_sc_hd__nand2_8 _18101_ (.A(_06002_),
    .B(_06711_),
    .Y(_06712_));
 sky130_fd_sc_hd__clkinv_8 _18102_ (.A(_06712_),
    .Y(\hash.CA1.S1.X[29] ));
 sky130_fd_sc_hd__a41oi_2 _18103_ (.A1(_06683_),
    .A2(_06684_),
    .A3(net1056),
    .A4(net1124),
    .B1(net1097),
    .Y(_06713_));
 sky130_fd_sc_hd__xnor2_2 _18104_ (.A(\hash.CA1.S1.X[29] ),
    .B(_06713_),
    .Y(_00802_));
 sky130_fd_sc_hd__nor4_2 _18105_ (.A(net345),
    .B(_13519_),
    .C(_13514_),
    .D(_13516_),
    .Y(_06714_));
 sky130_fd_sc_hd__nand3_1 _18106_ (.A(_06002_),
    .B(_13517_),
    .C(_13519_),
    .Y(_06715_));
 sky130_fd_sc_hd__nor2_4 _18107_ (.A(_06705_),
    .B(_06715_),
    .Y(_06716_));
 sky130_fd_sc_hd__nor4_1 _18108_ (.A(net345),
    .B(_13517_),
    .C(_13519_),
    .D(_13516_),
    .Y(_06717_));
 sky130_fd_sc_hd__a31oi_1 _18109_ (.A1(_06002_),
    .A2(_13519_),
    .A3(_13516_),
    .B1(_06717_),
    .Y(_06718_));
 sky130_fd_sc_hd__nand4_1 _18110_ (.A(_06002_),
    .B(_13517_),
    .C(_13519_),
    .D(_13514_),
    .Y(_06719_));
 sky130_fd_sc_hd__nand2_2 _18111_ (.A(_06718_),
    .B(_06719_),
    .Y(_06720_));
 sky130_fd_sc_hd__a211oi_4 _18112_ (.A1(_06705_),
    .A2(_06714_),
    .B1(_06720_),
    .C1(_06716_),
    .Y(\hash.CA1.S1.X[30] ));
 sky130_fd_sc_hd__a41o_1 _18113_ (.A1(_06674_),
    .A2(net1054),
    .A3(net1056),
    .A4(net1124),
    .B1(net1097),
    .X(_06721_));
 sky130_fd_sc_hd__nand2_2 _18114_ (.A(_06721_),
    .B(\hash.CA1.S1.X[29] ),
    .Y(_06722_));
 sky130_fd_sc_hd__xor2_2 _18115_ (.A(net1040),
    .B(_06722_),
    .X(_00804_));
 sky130_fd_sc_hd__nand2_1 _18116_ (.A(_13517_),
    .B(_13519_),
    .Y(_06723_));
 sky130_fd_sc_hd__a21oi_1 _18117_ (.A1(_13519_),
    .A2(_13516_),
    .B1(_13518_),
    .Y(_06724_));
 sky130_fd_sc_hd__o21ai_2 _18118_ (.A1(_06710_),
    .A2(_06723_),
    .B1(_06724_),
    .Y(_06725_));
 sky130_fd_sc_hd__xnor2_2 _18119_ (.A(\hash.CA2.p5[31] ),
    .B(_06248_),
    .Y(_06726_));
 sky130_fd_sc_hd__xnor2_2 _18120_ (.A(_06725_),
    .B(_06726_),
    .Y(_06727_));
 sky130_fd_sc_hd__nor2_4 _18121_ (.A(net534),
    .B(_06727_),
    .Y(\hash.CA1.S1.X[31] ));
 sky130_fd_sc_hd__o21ba_4 _18122_ (.A1(_06712_),
    .A2(_06713_),
    .B1_N(net1040),
    .X(_06728_));
 sky130_fd_sc_hd__xnor2_2 _18123_ (.A(\hash.CA1.S1.X[31] ),
    .B(_06728_),
    .Y(_00805_));
 sky130_fd_sc_hd__nand2_8 _18124_ (.A(_06002_),
    .B(\hash.CA2.b_dash[2] ),
    .Y(_12666_));
 sky130_fd_sc_hd__inv_1 _18125_ (.A(_12666_),
    .Y(_13857_));
 sky130_fd_sc_hd__nor2_4 _18126_ (.A(net343),
    .B(\hash.CA2.b_dash[3] ),
    .Y(_12674_));
 sky130_fd_sc_hd__xor2_1 _18127_ (.A(_13858_),
    .B(_12674_),
    .X(_00772_));
 sky130_fd_sc_hd__nor2_4 _18128_ (.A(net344),
    .B(\hash.CA2.b_dash[4] ),
    .Y(_12679_));
 sky130_fd_sc_hd__a21oi_1 _18129_ (.A1(\hash.CA2.b_dash[1] ),
    .A2(\hash.CA2.b_dash[2] ),
    .B1(\hash.CA2.b_dash[3] ),
    .Y(_06729_));
 sky130_fd_sc_hd__xnor2_1 _18130_ (.A(\hash.CA2.b_dash[4] ),
    .B(_06729_),
    .Y(_06730_));
 sky130_fd_sc_hd__nand2_1 _18131_ (.A(_06002_),
    .B(_06730_),
    .Y(_00774_));
 sky130_fd_sc_hd__or2_4 _18132_ (.A(net343),
    .B(\hash.CA2.b_dash[5] ),
    .X(_12684_));
 sky130_fd_sc_hd__nor4_1 _18133_ (.A(net343),
    .B(\hash.CA2.b_dash[3] ),
    .C(\hash.CA2.b_dash[4] ),
    .D(_13858_),
    .Y(_06731_));
 sky130_fd_sc_hd__xor2_1 _18134_ (.A(_12684_),
    .B(_06731_),
    .X(_00775_));
 sky130_fd_sc_hd__nand2b_4 _18135_ (.A_N(net340),
    .B(\hash.CA2.b_dash[6] ),
    .Y(_12692_));
 sky130_fd_sc_hd__nor3_1 _18136_ (.A(net343),
    .B(\hash.CA2.b_dash[3] ),
    .C(\hash.CA2.b_dash[4] ),
    .Y(_06732_));
 sky130_fd_sc_hd__a21oi_2 _18137_ (.A1(\hash.CA2.b_dash[1] ),
    .A2(\hash.CA2.b_dash[2] ),
    .B1(\hash.CA2.b_dash[5] ),
    .Y(_06733_));
 sky130_fd_sc_hd__nand2_1 _18138_ (.A(_06732_),
    .B(_06733_),
    .Y(_06734_));
 sky130_fd_sc_hd__xnor2_1 _18139_ (.A(_12692_),
    .B(_06734_),
    .Y(_00776_));
 sky130_fd_sc_hd__nor4_1 _18140_ (.A(\hash.CA2.b_dash[3] ),
    .B(\hash.CA2.b_dash[4] ),
    .C(\hash.CA2.b_dash[5] ),
    .D(_13858_),
    .Y(_06735_));
 sky130_fd_sc_hd__nor2_2 _18141_ (.A(_12692_),
    .B(_06735_),
    .Y(_06736_));
 sky130_fd_sc_hd__nand2_8 _18142_ (.A(_06002_),
    .B(\hash.CA2.b_dash[7] ),
    .Y(_12701_));
 sky130_fd_sc_hd__inv_1 _18143_ (.A(\hash.CA2.b_dash[7] ),
    .Y(_06737_));
 sky130_fd_sc_hd__nand2_1 _18144_ (.A(_06737_),
    .B(_06736_),
    .Y(_06738_));
 sky130_fd_sc_hd__o21ai_0 _18145_ (.A1(_06736_),
    .A2(_12701_),
    .B1(_06738_),
    .Y(_00777_));
 sky130_fd_sc_hd__nor2_4 _18146_ (.A(net344),
    .B(\hash.CA2.b_dash[8] ),
    .Y(_12708_));
 sky130_fd_sc_hd__a211oi_2 _18147_ (.A1(_06732_),
    .A2(_06733_),
    .B1(_12692_),
    .C1(_06737_),
    .Y(_06739_));
 sky130_fd_sc_hd__xor2_1 _18148_ (.A(_12708_),
    .B(_06739_),
    .X(_00778_));
 sky130_fd_sc_hd__clkinv_2 _18149_ (.A(\hash.CA2.b_dash[9] ),
    .Y(_06740_));
 sky130_fd_sc_hd__a21oi_2 _18150_ (.A1(\hash.CA2.b_dash[7] ),
    .A2(_06736_),
    .B1(\hash.CA2.b_dash[8] ),
    .Y(_06741_));
 sky130_fd_sc_hd__xnor2_1 _18151_ (.A(_06740_),
    .B(_06741_),
    .Y(_06742_));
 sky130_fd_sc_hd__nand2_1 _18152_ (.A(_06002_),
    .B(_06742_),
    .Y(_00779_));
 sky130_fd_sc_hd__nor2_4 _18153_ (.A(net344),
    .B(\hash.CA2.b_dash[10] ),
    .Y(_12723_));
 sky130_fd_sc_hd__nand2_8 _18154_ (.A(_06002_),
    .B(\hash.CA2.b_dash[9] ),
    .Y(_12714_));
 sky130_fd_sc_hd__nor2_1 _18155_ (.A(\hash.CA2.b_dash[8] ),
    .B(_06739_),
    .Y(_06743_));
 sky130_fd_sc_hd__nor2_1 _18156_ (.A(_12714_),
    .B(_06743_),
    .Y(_06744_));
 sky130_fd_sc_hd__mux2_1 _18157_ (.A0(_12723_),
    .A1(\hash.CA2.b_dash[10] ),
    .S(_06744_),
    .X(_00780_));
 sky130_fd_sc_hd__nand2_4 _18158_ (.A(_06002_),
    .B(\hash.CA2.b_dash[11] ),
    .Y(_06745_));
 sky130_fd_sc_hd__inv_8 _18159_ (.A(_06745_),
    .Y(_12732_));
 sky130_fd_sc_hd__o21ai_4 _18160_ (.A1(_06740_),
    .A2(_06741_),
    .B1(_12723_),
    .Y(_06746_));
 sky130_fd_sc_hd__xnor2_1 _18161_ (.A(_06745_),
    .B(_06746_),
    .Y(_00752_));
 sky130_fd_sc_hd__or2_4 _18162_ (.A(net344),
    .B(\hash.CA2.b_dash[12] ),
    .X(_06747_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1134 ();
 sky130_fd_sc_hd__inv_1 _18164_ (.A(\hash.CA2.b_dash[10] ),
    .Y(_06748_));
 sky130_fd_sc_hd__o21ai_0 _18165_ (.A1(\hash.CA2.b_dash[8] ),
    .A2(_06739_),
    .B1(\hash.CA2.b_dash[9] ),
    .Y(_06749_));
 sky130_fd_sc_hd__a21oi_2 _18166_ (.A1(_06748_),
    .A2(_06749_),
    .B1(_06745_),
    .Y(_06750_));
 sky130_fd_sc_hd__xnor2_1 _18167_ (.A(_06747_),
    .B(_06750_),
    .Y(_00753_));
 sky130_fd_sc_hd__nand2_1 _18168_ (.A(\hash.CA2.b_dash[7] ),
    .B(_06736_),
    .Y(_06751_));
 sky130_fd_sc_hd__a21oi_1 _18169_ (.A1(_12708_),
    .A2(_06751_),
    .B1(_12714_),
    .Y(_06752_));
 sky130_fd_sc_hd__o21a_4 _18170_ (.A1(\hash.CA2.b_dash[10] ),
    .A2(_06752_),
    .B1(\hash.CA2.b_dash[11] ),
    .X(_06753_));
 sky130_fd_sc_hd__nor2_1 _18171_ (.A(_06747_),
    .B(_06753_),
    .Y(_06754_));
 sky130_fd_sc_hd__or2_4 _18172_ (.A(net344),
    .B(\hash.CA2.b_dash[13] ),
    .X(_12746_));
 sky130_fd_sc_hd__nor2_1 _18173_ (.A(_06754_),
    .B(_12746_),
    .Y(_06755_));
 sky130_fd_sc_hd__a21oi_1 _18174_ (.A1(\hash.CA2.b_dash[13] ),
    .A2(_06754_),
    .B1(_06755_),
    .Y(_00754_));
 sky130_fd_sc_hd__nor2_4 _18175_ (.A(net345),
    .B(\hash.CA2.b_dash[14] ),
    .Y(_12752_));
 sky130_fd_sc_hd__o21ai_1 _18176_ (.A1(\hash.CA2.b_dash[10] ),
    .A2(_06744_),
    .B1(\hash.CA2.b_dash[11] ),
    .Y(_06756_));
 sky130_fd_sc_hd__nor2_1 _18177_ (.A(\hash.CA2.b_dash[13] ),
    .B(_06747_),
    .Y(_06757_));
 sky130_fd_sc_hd__nand2_2 _18178_ (.A(_06756_),
    .B(_06757_),
    .Y(_06758_));
 sky130_fd_sc_hd__xor2_1 _18179_ (.A(_12752_),
    .B(_06758_),
    .X(_00755_));
 sky130_fd_sc_hd__nor2_2 _18180_ (.A(net534),
    .B(\hash.CA2.b_dash[15] ),
    .Y(_12759_));
 sky130_fd_sc_hd__nor2_1 _18181_ (.A(\hash.CA2.b_dash[12] ),
    .B(\hash.CA2.b_dash[13] ),
    .Y(_06759_));
 sky130_fd_sc_hd__nand2_2 _18182_ (.A(_12752_),
    .B(_06759_),
    .Y(_06760_));
 sky130_fd_sc_hd__a21oi_4 _18183_ (.A1(_12732_),
    .A2(_06746_),
    .B1(_06760_),
    .Y(_06761_));
 sky130_fd_sc_hd__nor3_1 _18184_ (.A(net344),
    .B(\hash.CA2.b_dash[15] ),
    .C(_06761_),
    .Y(_06762_));
 sky130_fd_sc_hd__a21oi_1 _18185_ (.A1(\hash.CA2.b_dash[15] ),
    .A2(_06761_),
    .B1(_06762_),
    .Y(_00756_));
 sky130_fd_sc_hd__or2_4 _18186_ (.A(net344),
    .B(\hash.CA2.b_dash[16] ),
    .X(_12767_));
 sky130_fd_sc_hd__or2_4 _18187_ (.A(_06750_),
    .B(_06760_),
    .X(_06763_));
 sky130_fd_sc_hd__nor2_1 _18188_ (.A(\hash.CA2.b_dash[15] ),
    .B(_06763_),
    .Y(_06764_));
 sky130_fd_sc_hd__xor2_1 _18189_ (.A(_12767_),
    .B(_06764_),
    .X(_00757_));
 sky130_fd_sc_hd__nor2_4 _18190_ (.A(net344),
    .B(\hash.CA2.b_dash[17] ),
    .Y(_06765_));
 sky130_fd_sc_hd__inv_6 _18191_ (.A(_06765_),
    .Y(_12774_));
 sky130_fd_sc_hd__nor4_1 _18192_ (.A(net344),
    .B(\hash.CA2.b_dash[14] ),
    .C(\hash.CA2.b_dash[15] ),
    .D(\hash.CA2.b_dash[16] ),
    .Y(_06766_));
 sky130_fd_sc_hd__nand3b_1 _18193_ (.A_N(\hash.CA2.b_dash[13] ),
    .B(_06754_),
    .C(_06766_),
    .Y(_06767_));
 sky130_fd_sc_hd__xnor2_1 _18194_ (.A(_12774_),
    .B(_06767_),
    .Y(_00758_));
 sky130_fd_sc_hd__or2_4 _18195_ (.A(net343),
    .B(\hash.CA2.b_dash[18] ),
    .X(_12780_));
 sky130_fd_sc_hd__nor3b_1 _18196_ (.A(\hash.CA2.b_dash[17] ),
    .B(_06758_),
    .C_N(_06766_),
    .Y(_06768_));
 sky130_fd_sc_hd__xor2_1 _18197_ (.A(_12780_),
    .B(_06768_),
    .X(_00759_));
 sky130_fd_sc_hd__or2_4 _18198_ (.A(net344),
    .B(\hash.CA2.b_dash[19] ),
    .X(_12786_));
 sky130_fd_sc_hd__nor4_2 _18199_ (.A(net343),
    .B(\hash.CA2.b_dash[15] ),
    .C(\hash.CA2.b_dash[16] ),
    .D(\hash.CA2.b_dash[18] ),
    .Y(_06769_));
 sky130_fd_sc_hd__nand3_2 _18200_ (.A(_06761_),
    .B(_06765_),
    .C(_06769_),
    .Y(_06770_));
 sky130_fd_sc_hd__xnor2_1 _18201_ (.A(_12786_),
    .B(_06770_),
    .Y(_00760_));
 sky130_fd_sc_hd__nor2b_4 _18202_ (.A(net344),
    .B_N(\hash.CA2.b_dash[20] ),
    .Y(_06771_));
 sky130_fd_sc_hd__nor4b_4 _18203_ (.A(\hash.CA2.b_dash[17] ),
    .B(_06763_),
    .C(_12786_),
    .D_N(_06769_),
    .Y(_06772_));
 sky130_fd_sc_hd__xnor2_1 _18204_ (.A(_06771_),
    .B(_06772_),
    .Y(_00761_));
 sky130_fd_sc_hd__nor2b_1 _18205_ (.A(net534),
    .B_N(\hash.CA2.b_dash[21] ),
    .Y(_12802_));
 sky130_fd_sc_hd__o21a_4 _18206_ (.A1(\hash.CA2.b_dash[19] ),
    .A2(_06770_),
    .B1(\hash.CA2.b_dash[20] ),
    .X(_06773_));
 sky130_fd_sc_hd__xnor2_1 _18207_ (.A(\hash.CA2.b_dash[21] ),
    .B(_06773_),
    .Y(_06774_));
 sky130_fd_sc_hd__nor2_1 _18208_ (.A(net344),
    .B(_06774_),
    .Y(_00762_));
 sky130_fd_sc_hd__nor2_4 _18209_ (.A(net345),
    .B(\hash.CA2.b_dash[22] ),
    .Y(_12810_));
 sky130_fd_sc_hd__nand3b_1 _18210_ (.A_N(_06772_),
    .B(_06771_),
    .C(\hash.CA2.b_dash[21] ),
    .Y(_06775_));
 sky130_fd_sc_hd__xnor2_1 _18211_ (.A(_12810_),
    .B(_06775_),
    .Y(_00763_));
 sky130_fd_sc_hd__nor2b_4 _18212_ (.A(net345),
    .B_N(\hash.CA2.b_dash[23] ),
    .Y(_12818_));
 sky130_fd_sc_hd__a211o_4 _18213_ (.A1(\hash.CA2.b_dash[21] ),
    .A2(_06773_),
    .B1(\hash.CA2.b_dash[22] ),
    .C1(net345),
    .X(_06776_));
 sky130_fd_sc_hd__xor2_1 _18214_ (.A(_12818_),
    .B(_06776_),
    .X(_00764_));
 sky130_fd_sc_hd__nor2_4 _18215_ (.A(net345),
    .B(\hash.CA2.b_dash[24] ),
    .Y(_12826_));
 sky130_fd_sc_hd__nand2b_2 _18216_ (.A_N(\hash.CA2.b_dash[22] ),
    .B(_06775_),
    .Y(_06777_));
 sky130_fd_sc_hd__nand2_1 _18217_ (.A(_12818_),
    .B(_06777_),
    .Y(_06778_));
 sky130_fd_sc_hd__xnor2_1 _18218_ (.A(_12826_),
    .B(_06778_),
    .Y(_00765_));
 sky130_fd_sc_hd__nor2_4 _18219_ (.A(net342),
    .B(_04733_),
    .Y(_12834_));
 sky130_fd_sc_hd__a21boi_0 _18220_ (.A1(_12818_),
    .A2(_06776_),
    .B1_N(_12826_),
    .Y(_06779_));
 sky130_fd_sc_hd__xnor2_1 _18221_ (.A(_12834_),
    .B(_06779_),
    .Y(_00766_));
 sky130_fd_sc_hd__a21o_1 _18222_ (.A1(\hash.CA2.b_dash[23] ),
    .A2(_06777_),
    .B1(\hash.CA2.b_dash[24] ),
    .X(_06780_));
 sky130_fd_sc_hd__nand2_2 _18223_ (.A(_12834_),
    .B(_06780_),
    .Y(_06781_));
 sky130_fd_sc_hd__nor2_4 _18224_ (.A(net345),
    .B(\hash.CA2.b_dash[26] ),
    .Y(_06782_));
 sky130_fd_sc_hd__xnor2_1 _18225_ (.A(_06781_),
    .B(_06782_),
    .Y(_00767_));
 sky130_fd_sc_hd__nor2b_4 _18226_ (.A(net342),
    .B_N(\hash.CA2.b_dash[27] ),
    .Y(_12849_));
 sky130_fd_sc_hd__a21oi_1 _18227_ (.A1(\hash.CA2.b_dash[23] ),
    .A2(_06776_),
    .B1(\hash.CA2.b_dash[24] ),
    .Y(_06783_));
 sky130_fd_sc_hd__o21ai_2 _18228_ (.A1(_04733_),
    .A2(_06783_),
    .B1(_06782_),
    .Y(_06784_));
 sky130_fd_sc_hd__xor2_1 _18229_ (.A(_12849_),
    .B(_06784_),
    .X(_00768_));
 sky130_fd_sc_hd__inv_1 _18230_ (.A(\hash.CA2.b_dash[28] ),
    .Y(_06785_));
 sky130_fd_sc_hd__nor2_2 _18231_ (.A(net342),
    .B(_06785_),
    .Y(_12857_));
 sky130_fd_sc_hd__a21boi_2 _18232_ (.A1(_06781_),
    .A2(_06782_),
    .B1_N(_12849_),
    .Y(_06786_));
 sky130_fd_sc_hd__mux2_1 _18233_ (.A0(_12857_),
    .A1(_06785_),
    .S(_06786_),
    .X(_00769_));
 sky130_fd_sc_hd__or2_4 _18234_ (.A(net342),
    .B(\hash.CA2.b_dash[29] ),
    .X(_12864_));
 sky130_fd_sc_hd__and3_4 _18235_ (.A(\hash.CA2.b_dash[28] ),
    .B(_12849_),
    .C(_06784_),
    .X(_06787_));
 sky130_fd_sc_hd__xnor2_1 _18236_ (.A(_12864_),
    .B(_06787_),
    .Y(_00770_));
 sky130_fd_sc_hd__nor2b_2 _18237_ (.A(net534),
    .B_N(\hash.CA2.b_dash[30] ),
    .Y(_12871_));
 sky130_fd_sc_hd__a21oi_1 _18238_ (.A1(\hash.CA2.b_dash[28] ),
    .A2(_06786_),
    .B1(\hash.CA2.b_dash[29] ),
    .Y(_06788_));
 sky130_fd_sc_hd__xor2_1 _18239_ (.A(\hash.CA2.b_dash[30] ),
    .B(_06788_),
    .X(_06789_));
 sky130_fd_sc_hd__nand2_1 _18240_ (.A(_06002_),
    .B(_06789_),
    .Y(_00771_));
 sky130_fd_sc_hd__o21ai_0 _18241_ (.A1(\hash.CA2.b_dash[29] ),
    .A2(_06787_),
    .B1(\hash.CA2.b_dash[30] ),
    .Y(_06790_));
 sky130_fd_sc_hd__xnor2_1 _18242_ (.A(\hash.CA2.b_dash[31] ),
    .B(_06790_),
    .Y(_06791_));
 sky130_fd_sc_hd__nor2_1 _18243_ (.A(net342),
    .B(_06791_),
    .Y(_00773_));
 sky130_fd_sc_hd__xor2_1 _18244_ (.A(_13859_),
    .B(_13679_),
    .X(_00742_));
 sky130_fd_sc_hd__nand3_2 _18245_ (.A(\hash.CA2.a_dash[1] ),
    .B(\hash.CA2.a_dash[2] ),
    .C(\hash.CA2.a_dash[3] ),
    .Y(_06792_));
 sky130_fd_sc_hd__xnor2_1 _18246_ (.A(\hash.CA2.a_dash[4] ),
    .B(_06792_),
    .Y(_06793_));
 sky130_fd_sc_hd__nor2_1 _18247_ (.A(net340),
    .B(_06793_),
    .Y(_00744_));
 sky130_fd_sc_hd__or2_4 _18248_ (.A(net340),
    .B(\hash.CA2.a_dash[4] ),
    .X(_13685_));
 sky130_fd_sc_hd__a21oi_1 _18249_ (.A1(\hash.CA2.a_dash[3] ),
    .A2(_13859_),
    .B1(\hash.CA2.a_dash[4] ),
    .Y(_06794_));
 sky130_fd_sc_hd__xnor2_1 _18250_ (.A(\hash.CA2.a_dash[5] ),
    .B(_06794_),
    .Y(_06795_));
 sky130_fd_sc_hd__nand2_1 _18251_ (.A(_06002_),
    .B(_06795_),
    .Y(_00745_));
 sky130_fd_sc_hd__nor2_4 _18252_ (.A(\hash.CA2.a_dash[5] ),
    .B(_13685_),
    .Y(_06796_));
 sky130_fd_sc_hd__nand2_4 _18253_ (.A(_06792_),
    .B(_06796_),
    .Y(_06797_));
 sky130_fd_sc_hd__xnor2_1 _18254_ (.A(_13697_),
    .B(_06797_),
    .Y(_00746_));
 sky130_fd_sc_hd__a21oi_1 _18255_ (.A1(\hash.CA2.a_dash[3] ),
    .A2(_13859_),
    .B1(\hash.CA2.a_dash[6] ),
    .Y(_06798_));
 sky130_fd_sc_hd__nand2_4 _18256_ (.A(_06796_),
    .B(_06798_),
    .Y(_06799_));
 sky130_fd_sc_hd__nand2_8 _18257_ (.A(_06002_),
    .B(\hash.CA2.a_dash[7] ),
    .Y(_06800_));
 sky130_fd_sc_hd__xnor2_1 _18258_ (.A(_06799_),
    .B(_06800_),
    .Y(_00747_));
 sky130_fd_sc_hd__or2_0 _18259_ (.A(net346),
    .B(\hash.CA2.a_dash[8] ),
    .X(_13710_));
 sky130_fd_sc_hd__o21ai_0 _18260_ (.A1(\hash.CA2.a_dash[6] ),
    .A2(_06797_),
    .B1(\hash.CA2.a_dash[7] ),
    .Y(_06801_));
 sky130_fd_sc_hd__xnor2_1 _18261_ (.A(\hash.CA2.a_dash[8] ),
    .B(_06801_),
    .Y(_06802_));
 sky130_fd_sc_hd__nor2_1 _18262_ (.A(net340),
    .B(_06802_),
    .Y(_00748_));
 sky130_fd_sc_hd__a21oi_2 _18263_ (.A1(\hash.CA2.a_dash[7] ),
    .A2(_06799_),
    .B1(\hash.CA2.a_dash[8] ),
    .Y(_06803_));
 sky130_fd_sc_hd__xnor2_1 _18264_ (.A(\hash.CA2.a_dash[9] ),
    .B(_06803_),
    .Y(_06804_));
 sky130_fd_sc_hd__nand2_1 _18265_ (.A(_06002_),
    .B(_06804_),
    .Y(_00749_));
 sky130_fd_sc_hd__nor2b_4 _18266_ (.A(net340),
    .B_N(\hash.CA2.a_dash[10] ),
    .Y(_13721_));
 sky130_fd_sc_hd__nor2_2 _18267_ (.A(\hash.CA2.a_dash[6] ),
    .B(_06797_),
    .Y(_06805_));
 sky130_fd_sc_hd__nor2_1 _18268_ (.A(\hash.CA2.a_dash[8] ),
    .B(_13716_),
    .Y(_06806_));
 sky130_fd_sc_hd__o21ai_2 _18269_ (.A1(_06800_),
    .A2(_06805_),
    .B1(_06806_),
    .Y(_06807_));
 sky130_fd_sc_hd__xor2_1 _18270_ (.A(_13721_),
    .B(_06807_),
    .X(_00750_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1133 ();
 sky130_fd_sc_hd__clkinv_1 _18272_ (.A(_06803_),
    .Y(_06809_));
 sky130_fd_sc_hd__o21ai_0 _18273_ (.A1(\hash.CA2.a_dash[9] ),
    .A2(_06809_),
    .B1(\hash.CA2.a_dash[10] ),
    .Y(_06810_));
 sky130_fd_sc_hd__xor2_1 _18274_ (.A(\hash.CA2.a_dash[11] ),
    .B(_06810_),
    .X(_06811_));
 sky130_fd_sc_hd__nor2_1 _18275_ (.A(net340),
    .B(_06811_),
    .Y(_00722_));
 sky130_fd_sc_hd__or2_4 _18276_ (.A(net341),
    .B(\hash.CA2.a_dash[12] ),
    .X(_13734_));
 sky130_fd_sc_hd__and3_4 _18277_ (.A(\hash.CA2.a_dash[11] ),
    .B(_13721_),
    .C(_06807_),
    .X(_06812_));
 sky130_fd_sc_hd__xnor2_1 _18278_ (.A(_13734_),
    .B(_06812_),
    .Y(_00723_));
 sky130_fd_sc_hd__o211a_4 _18279_ (.A1(_13716_),
    .A2(_06809_),
    .B1(_13721_),
    .C1(\hash.CA2.a_dash[11] ),
    .X(_06813_));
 sky130_fd_sc_hd__or3_1 _18280_ (.A(\hash.CA2.a_dash[12] ),
    .B(\hash.CA2.a_dash[13] ),
    .C(_06813_),
    .X(_06814_));
 sky130_fd_sc_hd__o21ai_0 _18281_ (.A1(\hash.CA2.a_dash[12] ),
    .A2(_06813_),
    .B1(\hash.CA2.a_dash[13] ),
    .Y(_06815_));
 sky130_fd_sc_hd__nand3_1 _18282_ (.A(_06002_),
    .B(_06814_),
    .C(_06815_),
    .Y(_00724_));
 sky130_fd_sc_hd__or3_4 _18283_ (.A(net341),
    .B(\hash.CA2.a_dash[12] ),
    .C(\hash.CA2.a_dash[13] ),
    .X(_06816_));
 sky130_fd_sc_hd__nor2_1 _18284_ (.A(_06812_),
    .B(_06816_),
    .Y(_06817_));
 sky130_fd_sc_hd__xor2_1 _18285_ (.A(_13746_),
    .B(_06817_),
    .X(_00725_));
 sky130_fd_sc_hd__or3_4 _18286_ (.A(\hash.CA2.a_dash[14] ),
    .B(_06813_),
    .C(_06816_),
    .X(_06818_));
 sky130_fd_sc_hd__xnor2_1 _18287_ (.A(_13753_),
    .B(_06818_),
    .Y(_00726_));
 sky130_fd_sc_hd__nor2b_4 _18288_ (.A(net341),
    .B_N(\hash.CA2.a_dash[16] ),
    .Y(_13760_));
 sky130_fd_sc_hd__or4_4 _18289_ (.A(\hash.CA2.a_dash[15] ),
    .B(_13746_),
    .C(_06812_),
    .D(_06816_),
    .X(_06819_));
 sky130_fd_sc_hd__xor2_1 _18290_ (.A(_13760_),
    .B(_06819_),
    .X(_00727_));
 sky130_fd_sc_hd__nor2_2 _18291_ (.A(net341),
    .B(\hash.CA2.a_dash[17] ),
    .Y(_06820_));
 sky130_fd_sc_hd__inv_4 _18292_ (.A(_06820_),
    .Y(_13767_));
 sky130_fd_sc_hd__o21ai_4 _18293_ (.A1(\hash.CA2.a_dash[15] ),
    .A2(_06818_),
    .B1(_13760_),
    .Y(_06821_));
 sky130_fd_sc_hd__mux2_1 _18294_ (.A0(\hash.CA2.a_dash[17] ),
    .A1(_06820_),
    .S(_06821_),
    .X(_00728_));
 sky130_fd_sc_hd__or2_0 _18295_ (.A(net346),
    .B(\hash.CA2.a_dash[18] ),
    .X(_13773_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1132 ();
 sky130_fd_sc_hd__a21oi_1 _18297_ (.A1(\hash.CA2.a_dash[16] ),
    .A2(_06819_),
    .B1(\hash.CA2.a_dash[17] ),
    .Y(_06823_));
 sky130_fd_sc_hd__xnor2_1 _18298_ (.A(\hash.CA2.a_dash[18] ),
    .B(_06823_),
    .Y(_06824_));
 sky130_fd_sc_hd__nand2_1 _18299_ (.A(_06002_),
    .B(_06824_),
    .Y(_00729_));
 sky130_fd_sc_hd__nand3b_1 _18300_ (.A_N(\hash.CA2.a_dash[18] ),
    .B(_06820_),
    .C(_06821_),
    .Y(_06825_));
 sky130_fd_sc_hd__xnor2_1 _18301_ (.A(_13778_),
    .B(_06825_),
    .Y(_00730_));
 sky130_fd_sc_hd__nor2b_4 _18302_ (.A(net341),
    .B_N(\hash.CA2.a_dash[20] ),
    .Y(_13783_));
 sky130_fd_sc_hd__nand2_1 _18303_ (.A(\hash.CA2.a_dash[16] ),
    .B(_06819_),
    .Y(_06826_));
 sky130_fd_sc_hd__nor3_2 _18304_ (.A(\hash.CA2.a_dash[18] ),
    .B(\hash.CA2.a_dash[19] ),
    .C(_13767_),
    .Y(_06827_));
 sky130_fd_sc_hd__nand2_2 _18305_ (.A(_06826_),
    .B(_06827_),
    .Y(_06828_));
 sky130_fd_sc_hd__xor2_1 _18306_ (.A(_13783_),
    .B(_06828_),
    .X(_00731_));
 sky130_fd_sc_hd__or2_4 _18307_ (.A(net346),
    .B(\hash.CA2.a_dash[21] ),
    .X(_13788_));
 sky130_fd_sc_hd__a21boi_4 _18308_ (.A1(_06821_),
    .A2(_06827_),
    .B1_N(\hash.CA2.a_dash[20] ),
    .Y(_06829_));
 sky130_fd_sc_hd__xor2_1 _18309_ (.A(\hash.CA2.a_dash[21] ),
    .B(_06829_),
    .X(_06830_));
 sky130_fd_sc_hd__nor2_1 _18310_ (.A(net343),
    .B(_06830_),
    .Y(_00732_));
 sky130_fd_sc_hd__or2_4 _18311_ (.A(net343),
    .B(\hash.CA2.a_dash[22] ),
    .X(_13793_));
 sky130_fd_sc_hd__a21oi_2 _18312_ (.A1(\hash.CA2.a_dash[20] ),
    .A2(_06828_),
    .B1(\hash.CA2.a_dash[21] ),
    .Y(_06831_));
 sky130_fd_sc_hd__xnor2_1 _18313_ (.A(\hash.CA2.a_dash[22] ),
    .B(_06831_),
    .Y(_06832_));
 sky130_fd_sc_hd__nand2_1 _18314_ (.A(_06002_),
    .B(_06832_),
    .Y(_00733_));
 sky130_fd_sc_hd__nor2b_4 _18315_ (.A(net343),
    .B_N(\hash.CA2.a_dash[23] ),
    .Y(_13799_));
 sky130_fd_sc_hd__or3_4 _18316_ (.A(\hash.CA2.a_dash[21] ),
    .B(_06829_),
    .C(_13793_),
    .X(_06833_));
 sky130_fd_sc_hd__xor2_1 _18317_ (.A(_13799_),
    .B(_06833_),
    .X(_00734_));
 sky130_fd_sc_hd__nand2b_1 _18318_ (.A_N(_13793_),
    .B(_06831_),
    .Y(_06834_));
 sky130_fd_sc_hd__nand2_1 _18319_ (.A(\hash.CA2.a_dash[23] ),
    .B(_06834_),
    .Y(_06835_));
 sky130_fd_sc_hd__xor2_1 _18320_ (.A(\hash.CA2.a_dash[24] ),
    .B(_06835_),
    .X(_06836_));
 sky130_fd_sc_hd__nor2_1 _18321_ (.A(net343),
    .B(_06836_),
    .Y(_00735_));
 sky130_fd_sc_hd__nand3_1 _18322_ (.A(\hash.CA2.a_dash[23] ),
    .B(\hash.CA2.a_dash[24] ),
    .C(_06833_),
    .Y(_06837_));
 sky130_fd_sc_hd__xnor2_1 _18323_ (.A(_04734_),
    .B(_06837_),
    .Y(_06838_));
 sky130_fd_sc_hd__nor2_1 _18324_ (.A(net343),
    .B(_06838_),
    .Y(_00736_));
 sky130_fd_sc_hd__nand4_1 _18325_ (.A(\hash.CA2.a_dash[24] ),
    .B(\hash.CA2.a_dash[25] ),
    .C(_13799_),
    .D(_06834_),
    .Y(_06839_));
 sky130_fd_sc_hd__xor2_1 _18326_ (.A(_06287_),
    .B(_06839_),
    .X(_00737_));
 sky130_fd_sc_hd__and4_4 _18327_ (.A(\hash.CA2.a_dash[24] ),
    .B(\hash.CA2.a_dash[25] ),
    .C(_13799_),
    .D(_06833_),
    .X(_06840_));
 sky130_fd_sc_hd__or3_1 _18328_ (.A(\hash.CA2.a_dash[26] ),
    .B(\hash.CA2.a_dash[27] ),
    .C(_06840_),
    .X(_06841_));
 sky130_fd_sc_hd__o21ai_0 _18329_ (.A1(\hash.CA2.a_dash[26] ),
    .A2(_06840_),
    .B1(\hash.CA2.a_dash[27] ),
    .Y(_06842_));
 sky130_fd_sc_hd__nand3_1 _18330_ (.A(_06002_),
    .B(_06841_),
    .C(_06842_),
    .Y(_00738_));
 sky130_fd_sc_hd__nor2_1 _18331_ (.A(\hash.CA2.a_dash[27] ),
    .B(_06287_),
    .Y(_06843_));
 sky130_fd_sc_hd__nand2_1 _18332_ (.A(_06839_),
    .B(_06843_),
    .Y(_06844_));
 sky130_fd_sc_hd__xnor2_1 _18333_ (.A(_13834_),
    .B(_06844_),
    .Y(_00739_));
 sky130_fd_sc_hd__or3_4 _18334_ (.A(\hash.CA2.a_dash[27] ),
    .B(\hash.CA2.a_dash[28] ),
    .C(_06287_),
    .X(_06845_));
 sky130_fd_sc_hd__nor2_1 _18335_ (.A(_06840_),
    .B(_06845_),
    .Y(_06846_));
 sky130_fd_sc_hd__xor2_1 _18336_ (.A(_13840_),
    .B(_06846_),
    .X(_00740_));
 sky130_fd_sc_hd__nor2_4 _18337_ (.A(net346),
    .B(_04769_),
    .Y(_13845_));
 sky130_fd_sc_hd__nor2_1 _18338_ (.A(\hash.CA2.a_dash[29] ),
    .B(_06845_),
    .Y(_06847_));
 sky130_fd_sc_hd__nand2_1 _18339_ (.A(_06839_),
    .B(_06847_),
    .Y(_06848_));
 sky130_fd_sc_hd__xor2_1 _18340_ (.A(_13845_),
    .B(_06848_),
    .X(_00741_));
 sky130_fd_sc_hd__o31ai_1 _18341_ (.A1(\hash.CA2.a_dash[29] ),
    .A2(_06840_),
    .A3(_06845_),
    .B1(\hash.CA2.a_dash[30] ),
    .Y(_06849_));
 sky130_fd_sc_hd__xor2_1 _18342_ (.A(\hash.CA2.a_dash[31] ),
    .B(_06849_),
    .X(_06850_));
 sky130_fd_sc_hd__nor2_1 _18343_ (.A(net343),
    .B(_06850_),
    .Y(_00743_));
 sky130_fd_sc_hd__xnor2_1 _18344_ (.A(_13860_),
    .B(\hash.CA1.b[2] ),
    .Y(_00711_));
 sky130_fd_sc_hd__a21oi_1 _18345_ (.A1(_12922_),
    .A2(_12082_),
    .B1(_04421_),
    .Y(_06851_));
 sky130_fd_sc_hd__xor2_1 _18346_ (.A(_04470_),
    .B(_06851_),
    .X(_06852_));
 sky130_fd_sc_hd__nand2_1 _18347_ (.A(_06002_),
    .B(_06852_),
    .Y(_00714_));
 sky130_fd_sc_hd__o21ai_0 _18348_ (.A1(_13860_),
    .A2(_04421_),
    .B1(_04470_),
    .Y(_06853_));
 sky130_fd_sc_hd__xor2_1 _18349_ (.A(_04487_),
    .B(_06853_),
    .X(_06854_));
 sky130_fd_sc_hd__nor2_1 _18350_ (.A(net340),
    .B(_06854_),
    .Y(_00715_));
 sky130_fd_sc_hd__and4bb_4 _18351_ (.A_N(net340),
    .B_N(_06851_),
    .C(_04487_),
    .D(_04470_),
    .X(_06855_));
 sky130_fd_sc_hd__xor2_1 _18352_ (.A(\hash.CA1.b[5] ),
    .B(_06855_),
    .X(_00716_));
 sky130_fd_sc_hd__o211a_4 _18353_ (.A1(_13860_),
    .A2(_04421_),
    .B1(_04470_),
    .C1(_04501_),
    .X(_06856_));
 sky130_fd_sc_hd__nand2_1 _18354_ (.A(\hash.CA1.b[4] ),
    .B(_06856_),
    .Y(_06857_));
 sky130_fd_sc_hd__xnor2_1 _18355_ (.A(\hash.CA1.b[6] ),
    .B(_06857_),
    .Y(_00717_));
 sky130_fd_sc_hd__nand3_1 _18356_ (.A(_04501_),
    .B(_04522_),
    .C(_06855_),
    .Y(_06858_));
 sky130_fd_sc_hd__xor2_1 _18357_ (.A(\hash.CA1.b[7] ),
    .B(_06858_),
    .X(_00718_));
 sky130_fd_sc_hd__xnor2_1 _18358_ (.A(_12930_),
    .B(_04400_),
    .Y(_06859_));
 sky130_fd_sc_hd__nand3_1 _18359_ (.A(_04487_),
    .B(_06856_),
    .C(_06859_),
    .Y(_06860_));
 sky130_fd_sc_hd__nand3_2 _18360_ (.A(_06002_),
    .B(_04543_),
    .C(_06860_),
    .Y(_06861_));
 sky130_fd_sc_hd__nor2_1 _18361_ (.A(_04562_),
    .B(_06861_),
    .Y(_06862_));
 sky130_fd_sc_hd__a21oi_1 _18362_ (.A1(_06279_),
    .A2(_06861_),
    .B1(_06862_),
    .Y(_00719_));
 sky130_fd_sc_hd__a31o_1 _18363_ (.A1(_04501_),
    .A2(_04522_),
    .A3(_06855_),
    .B1(_04542_),
    .X(_06863_));
 sky130_fd_sc_hd__and2_4 _18364_ (.A(_06279_),
    .B(_06863_),
    .X(_06864_));
 sky130_fd_sc_hd__nand2_1 _18365_ (.A(_04580_),
    .B(_06864_),
    .Y(_06865_));
 sky130_fd_sc_hd__o21ai_0 _18366_ (.A1(_06280_),
    .A2(_06864_),
    .B1(_06865_),
    .Y(_00720_));
 sky130_fd_sc_hd__nand3_1 _18367_ (.A(\hash.CA1.b[4] ),
    .B(\hash.CA1.b[6] ),
    .C(_06856_),
    .Y(_06866_));
 sky130_fd_sc_hd__nand2_1 _18368_ (.A(_04543_),
    .B(_06866_),
    .Y(_06867_));
 sky130_fd_sc_hd__a21oi_1 _18369_ (.A1(_04562_),
    .A2(_06867_),
    .B1(_04580_),
    .Y(_06868_));
 sky130_fd_sc_hd__xnor2_1 _18370_ (.A(_04599_),
    .B(_06868_),
    .Y(_06869_));
 sky130_fd_sc_hd__nand2_1 _18371_ (.A(_06002_),
    .B(_06869_),
    .Y(_00691_));
 sky130_fd_sc_hd__nor3_1 _18372_ (.A(_04580_),
    .B(\hash.CA1.b[10] ),
    .C(_06864_),
    .Y(_06870_));
 sky130_fd_sc_hd__xnor2_1 _18373_ (.A(_06282_),
    .B(_06870_),
    .Y(_00692_));
 sky130_fd_sc_hd__a2111o_2 _18374_ (.A1(_04562_),
    .A2(_06861_),
    .B1(_06280_),
    .C1(_04614_),
    .D1(_04599_),
    .X(_06871_));
 sky130_fd_sc_hd__xor2_1 _18375_ (.A(_06283_),
    .B(_06871_),
    .X(_00693_));
 sky130_fd_sc_hd__a2111o_2 _18376_ (.A1(_06279_),
    .A2(_06863_),
    .B1(_06280_),
    .C1(_04599_),
    .D1(_04614_),
    .X(_06872_));
 sky130_fd_sc_hd__nand2_1 _18377_ (.A(_04623_),
    .B(_06872_),
    .Y(_06873_));
 sky130_fd_sc_hd__xnor2_1 _18378_ (.A(_04437_),
    .B(_06873_),
    .Y(_06874_));
 sky130_fd_sc_hd__nor2_1 _18379_ (.A(net341),
    .B(_06874_),
    .Y(_00694_));
 sky130_fd_sc_hd__a21oi_2 _18380_ (.A1(_04623_),
    .A2(_06871_),
    .B1(_04437_),
    .Y(_06875_));
 sky130_fd_sc_hd__xnor2_1 _18381_ (.A(net1048),
    .B(_06875_),
    .Y(_06876_));
 sky130_fd_sc_hd__nand2_1 _18382_ (.A(_06002_),
    .B(_06876_),
    .Y(_00695_));
 sky130_fd_sc_hd__a21oi_4 _18383_ (.A1(_06283_),
    .A2(_06872_),
    .B1(_04437_),
    .Y(_06877_));
 sky130_fd_sc_hd__nor3_1 _18384_ (.A(net1046),
    .B(_04484_),
    .C(_06877_),
    .Y(_06878_));
 sky130_fd_sc_hd__o21a_1 _18385_ (.A1(net1046),
    .A2(_06877_),
    .B1(_04484_),
    .X(_06879_));
 sky130_fd_sc_hd__nor3_1 _18386_ (.A(net341),
    .B(_06878_),
    .C(_06879_),
    .Y(_00696_));
 sky130_fd_sc_hd__a21oi_1 _18387_ (.A1(_06283_),
    .A2(_06871_),
    .B1(_04437_),
    .Y(_06880_));
 sky130_fd_sc_hd__nor2_1 _18388_ (.A(net1047),
    .B(_06880_),
    .Y(_06881_));
 sky130_fd_sc_hd__nor2_1 _18389_ (.A(_04484_),
    .B(_06881_),
    .Y(_06882_));
 sky130_fd_sc_hd__xnor2_1 _18390_ (.A(_04503_),
    .B(_06882_),
    .Y(_06883_));
 sky130_fd_sc_hd__nand2_1 _18391_ (.A(_06002_),
    .B(_06883_),
    .Y(_00697_));
 sky130_fd_sc_hd__nor3_2 _18392_ (.A(net341),
    .B(_04484_),
    .C(_04503_),
    .Y(_06884_));
 sky130_fd_sc_hd__o21ai_4 _18393_ (.A1(net1044),
    .A2(_06877_),
    .B1(_06884_),
    .Y(_06885_));
 sky130_fd_sc_hd__xnor2_1 _18394_ (.A(\hash.CA1.b[17] ),
    .B(_06885_),
    .Y(_00698_));
 sky130_fd_sc_hd__o21ai_2 _18395_ (.A1(net1045),
    .A2(_06875_),
    .B1(_06884_),
    .Y(_06886_));
 sky130_fd_sc_hd__or2_4 _18396_ (.A(_04520_),
    .B(_06886_),
    .X(_06887_));
 sky130_fd_sc_hd__xnor2_1 _18397_ (.A(\hash.CA1.b[18] ),
    .B(_06887_),
    .Y(_00699_));
 sky130_fd_sc_hd__nor4_4 _18398_ (.A(net341),
    .B(_04520_),
    .C(_04541_),
    .D(_06885_),
    .Y(_06888_));
 sky130_fd_sc_hd__xnor2_1 _18399_ (.A(_06284_),
    .B(_06888_),
    .Y(_00700_));
 sky130_fd_sc_hd__o21ai_0 _18400_ (.A1(_04541_),
    .A2(_06887_),
    .B1(_04559_),
    .Y(_06889_));
 sky130_fd_sc_hd__xnor2_1 _18401_ (.A(_04681_),
    .B(_06889_),
    .Y(_06890_));
 sky130_fd_sc_hd__nor2_1 _18402_ (.A(net343),
    .B(_06890_),
    .Y(_00701_));
 sky130_fd_sc_hd__nand2_2 _18403_ (.A(_04577_),
    .B(_06284_),
    .Y(_06891_));
 sky130_fd_sc_hd__nor2_1 _18404_ (.A(_06888_),
    .B(_06891_),
    .Y(_06892_));
 sky130_fd_sc_hd__xnor2_1 _18405_ (.A(\hash.CA1.b[21] ),
    .B(_06892_),
    .Y(_00702_));
 sky130_fd_sc_hd__o311a_4 _18406_ (.A1(_04520_),
    .A2(_04541_),
    .A3(_06886_),
    .B1(_06284_),
    .C1(_04577_),
    .X(_06893_));
 sky130_fd_sc_hd__nor2_1 _18407_ (.A(\hash.CA1.b[21] ),
    .B(_06893_),
    .Y(_06894_));
 sky130_fd_sc_hd__xor2_1 _18408_ (.A(\hash.CA1.b[22] ),
    .B(_06894_),
    .X(_00703_));
 sky130_fd_sc_hd__clkinv_1 _18409_ (.A(_06285_),
    .Y(_06895_));
 sky130_fd_sc_hd__o21ai_2 _18410_ (.A1(_04420_),
    .A2(\hash.CA1.b[21] ),
    .B1(_06285_),
    .Y(_06896_));
 sky130_fd_sc_hd__o31ai_2 _18411_ (.A1(_06895_),
    .A2(_06888_),
    .A3(_06891_),
    .B1(_06896_),
    .Y(_06897_));
 sky130_fd_sc_hd__or3_1 _18412_ (.A(_04420_),
    .B(\hash.CA1.b[21] ),
    .C(_06892_),
    .X(_06898_));
 sky130_fd_sc_hd__nor2_1 _18413_ (.A(_06285_),
    .B(_06898_),
    .Y(_06899_));
 sky130_fd_sc_hd__nor2_1 _18414_ (.A(_06897_),
    .B(_06899_),
    .Y(_00704_));
 sky130_fd_sc_hd__o31ai_1 _18415_ (.A1(_04420_),
    .A2(\hash.CA1.b[21] ),
    .A3(_06893_),
    .B1(_04467_),
    .Y(_06900_));
 sky130_fd_sc_hd__xnor2_1 _18416_ (.A(_04726_),
    .B(_06900_),
    .Y(_06901_));
 sky130_fd_sc_hd__nor2_1 _18417_ (.A(net343),
    .B(_06901_),
    .Y(_00705_));
 sky130_fd_sc_hd__a21oi_1 _18418_ (.A1(_04467_),
    .A2(_06898_),
    .B1(\hash.CA1.b[24] ),
    .Y(_06902_));
 sky130_fd_sc_hd__xor2_1 _18419_ (.A(\hash.CA1.b[25] ),
    .B(_06902_),
    .X(_00706_));
 sky130_fd_sc_hd__nand2_1 _18420_ (.A(_06285_),
    .B(_06893_),
    .Y(_06903_));
 sky130_fd_sc_hd__nor2_1 _18421_ (.A(_04726_),
    .B(\hash.CA1.b[25] ),
    .Y(_06904_));
 sky130_fd_sc_hd__nand3_1 _18422_ (.A(_06896_),
    .B(_06903_),
    .C(_06904_),
    .Y(_06905_));
 sky130_fd_sc_hd__xor2_1 _18423_ (.A(\hash.CA1.b[26] ),
    .B(_06905_),
    .X(_00707_));
 sky130_fd_sc_hd__a21oi_1 _18424_ (.A1(_04481_),
    .A2(_04499_),
    .B1(net341),
    .Y(_06906_));
 sky130_fd_sc_hd__o21ai_2 _18425_ (.A1(_06897_),
    .A2(_06906_),
    .B1(net1102),
    .Y(_06907_));
 sky130_fd_sc_hd__xnor2_1 _18426_ (.A(_06288_),
    .B(_06907_),
    .Y(_00708_));
 sky130_fd_sc_hd__a31oi_2 _18427_ (.A1(_06896_),
    .A2(_06903_),
    .A3(_06904_),
    .B1(_06286_),
    .Y(_06908_));
 sky130_fd_sc_hd__or3_1 _18428_ (.A(net1070),
    .B(_04554_),
    .C(_06908_),
    .X(_06909_));
 sky130_fd_sc_hd__o21ai_0 _18429_ (.A1(net1069),
    .A2(_06908_),
    .B1(_04554_),
    .Y(_06910_));
 sky130_fd_sc_hd__nand3_1 _18430_ (.A(_06002_),
    .B(_06909_),
    .C(_06910_),
    .Y(_00709_));
 sky130_fd_sc_hd__nand2_1 _18431_ (.A(_06002_),
    .B(_04574_),
    .Y(\hash.CA1.b[29] ));
 sky130_fd_sc_hd__nor3b_1 _18432_ (.A(net1071),
    .B(_04554_),
    .C_N(_06907_),
    .Y(_06911_));
 sky130_fd_sc_hd__xnor2_1 _18433_ (.A(_04754_),
    .B(_06911_),
    .Y(_06912_));
 sky130_fd_sc_hd__nand2_1 _18434_ (.A(_06002_),
    .B(_06912_),
    .Y(_00710_));
 sky130_fd_sc_hd__nor4_1 _18435_ (.A(_04554_),
    .B(_04754_),
    .C(\hash.CA1.b[27] ),
    .D(_06908_),
    .Y(_06913_));
 sky130_fd_sc_hd__xnor2_1 _18436_ (.A(\hash.CA1.b[30] ),
    .B(_06913_),
    .Y(_00712_));
 sky130_fd_sc_hd__a41oi_1 _18437_ (.A1(_04662_),
    .A2(_04574_),
    .A3(_06288_),
    .A4(_06907_),
    .B1(_04588_),
    .Y(_06914_));
 sky130_fd_sc_hd__xor2_1 _18438_ (.A(net1078),
    .B(_06914_),
    .X(_06915_));
 sky130_fd_sc_hd__nor2_1 _18439_ (.A(net343),
    .B(_06915_),
    .Y(_00713_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1131 ();
 sky130_fd_sc_hd__nor2b_1 _18441_ (.A(net344),
    .B_N(\hash.CA2.S1.X[0] ),
    .Y(\hash.CA1.f[0] ));
 sky130_fd_sc_hd__mux2i_1 _18442_ (.A0(\hash.CA2.e_dash[0] ),
    .A1(\hash.CA2.S1.X[0] ),
    .S(_13445_),
    .Y(_06917_));
 sky130_fd_sc_hd__nor2_4 _18443_ (.A(net344),
    .B(_06917_),
    .Y(_13862_));
 sky130_fd_sc_hd__nor2b_1 _18444_ (.A(net344),
    .B_N(net1105),
    .Y(\hash.CA1.f[1] ));
 sky130_fd_sc_hd__mux2i_2 _18445_ (.A0(\hash.CA2.e_dash[1] ),
    .A1(\hash.CA2.S1.X[1] ),
    .S(_12365_),
    .Y(_06918_));
 sky130_fd_sc_hd__nor2_2 _18446_ (.A(net344),
    .B(_06918_),
    .Y(_12502_));
 sky130_fd_sc_hd__xor2_2 _18447_ (.A(_12498_),
    .B(_13868_),
    .X(_12509_));
 sky130_fd_sc_hd__inv_1 _18448_ (.A(_12509_),
    .Y(_12665_));
 sky130_fd_sc_hd__xor2_1 _18449_ (.A(_12503_),
    .B(_13872_),
    .X(_12508_));
 sky130_fd_sc_hd__inv_1 _18450_ (.A(_12508_),
    .Y(_12671_));
 sky130_fd_sc_hd__a21oi_4 _18451_ (.A1(_12497_),
    .A2(_13864_),
    .B1(_13863_),
    .Y(_06919_));
 sky130_fd_sc_hd__nor2b_1 _18452_ (.A(_06919_),
    .B_N(_13868_),
    .Y(_06920_));
 sky130_fd_sc_hd__nor2_1 _18453_ (.A(_13867_),
    .B(_06920_),
    .Y(_06921_));
 sky130_fd_sc_hd__xor2_2 _18454_ (.A(_13876_),
    .B(_06921_),
    .X(_12514_));
 sky130_fd_sc_hd__inv_1 _18455_ (.A(_13851_),
    .Y(\hash.CA1.f[3] ));
 sky130_fd_sc_hd__nor2_1 _18456_ (.A(\hash.CA2.e_dash[3] ),
    .B(\hash.CA1.S1.X[3] ),
    .Y(_06922_));
 sky130_fd_sc_hd__a21oi_4 _18457_ (.A1(_13851_),
    .A2(\hash.CA1.S1.X[3] ),
    .B1(_06922_),
    .Y(_13878_));
 sky130_fd_sc_hd__a21oi_2 _18458_ (.A1(_12500_),
    .A2(_13866_),
    .B1(_13865_),
    .Y(_06923_));
 sky130_fd_sc_hd__nor2b_4 _18459_ (.A(_06923_),
    .B_N(_13872_),
    .Y(_06924_));
 sky130_fd_sc_hd__nor2_1 _18460_ (.A(_13871_),
    .B(_06924_),
    .Y(_06925_));
 sky130_fd_sc_hd__xor2_2 _18461_ (.A(_13880_),
    .B(_06925_),
    .X(_12513_));
 sky130_fd_sc_hd__inv_2 _18462_ (.A(_13885_),
    .Y(_06926_));
 sky130_fd_sc_hd__a21o_1 _18463_ (.A1(_12498_),
    .A2(_13868_),
    .B1(_13867_),
    .X(_06927_));
 sky130_fd_sc_hd__a21oi_2 _18464_ (.A1(_13876_),
    .A2(_06927_),
    .B1(_13875_),
    .Y(_06928_));
 sky130_fd_sc_hd__xnor2_2 _18465_ (.A(_06926_),
    .B(_06928_),
    .Y(_12519_));
 sky130_fd_sc_hd__clkinvlp_4 _18466_ (.A(_13889_),
    .Y(_06929_));
 sky130_fd_sc_hd__a21o_1 _18467_ (.A1(_13872_),
    .A2(_12503_),
    .B1(_13871_),
    .X(_06930_));
 sky130_fd_sc_hd__a21oi_4 _18468_ (.A1(_13880_),
    .A2(_06930_),
    .B1(_13879_),
    .Y(_06931_));
 sky130_fd_sc_hd__xnor2_2 _18469_ (.A(_06929_),
    .B(_06931_),
    .Y(_12518_));
 sky130_fd_sc_hd__a21oi_1 _18470_ (.A1(_13880_),
    .A2(_13871_),
    .B1(_13879_),
    .Y(_06932_));
 sky130_fd_sc_hd__nor2_2 _18471_ (.A(_06929_),
    .B(_06932_),
    .Y(_06933_));
 sky130_fd_sc_hd__a311oi_1 _18472_ (.A1(_13880_),
    .A2(_13889_),
    .A3(_06924_),
    .B1(_06933_),
    .C1(_13888_),
    .Y(_06934_));
 sky130_fd_sc_hd__xnor2_1 _18473_ (.A(_13899_),
    .B(_06934_),
    .Y(_12523_));
 sky130_fd_sc_hd__inv_1 _18474_ (.A(_12523_),
    .Y(_12688_));
 sky130_fd_sc_hd__o21bai_2 _18475_ (.A1(_06926_),
    .A2(_06928_),
    .B1_N(_13884_),
    .Y(_06935_));
 sky130_fd_sc_hd__a21oi_4 _18476_ (.A1(_13895_),
    .A2(_06935_),
    .B1(_13894_),
    .Y(_06936_));
 sky130_fd_sc_hd__xnor2_2 _18477_ (.A(_13904_),
    .B(_06936_),
    .Y(_12529_));
 sky130_fd_sc_hd__inv_1 _18478_ (.A(_12529_),
    .Y(_12691_));
 sky130_fd_sc_hd__mux2_8 _18479_ (.A0(\hash.CA2.e_dash[6] ),
    .A1(\hash.CA1.f[6] ),
    .S(\hash.CA1.S1.X[6] ),
    .X(_13906_));
 sky130_fd_sc_hd__o21bai_1 _18480_ (.A1(_06931_),
    .A2(_06929_),
    .B1_N(_13888_),
    .Y(_06937_));
 sky130_fd_sc_hd__a21oi_2 _18481_ (.A1(_13899_),
    .A2(_06937_),
    .B1(_13898_),
    .Y(_06938_));
 sky130_fd_sc_hd__xnor2_1 _18482_ (.A(_13908_),
    .B(_06938_),
    .Y(_12528_));
 sky130_fd_sc_hd__inv_1 _18483_ (.A(_12528_),
    .Y(_12697_));
 sky130_fd_sc_hd__o21ai_0 _18484_ (.A1(_13895_),
    .A2(_13894_),
    .B1(_13904_),
    .Y(_06939_));
 sky130_fd_sc_hd__nand2b_2 _18485_ (.A_N(_13903_),
    .B(_06939_),
    .Y(_06940_));
 sky130_fd_sc_hd__a21o_1 _18486_ (.A1(_13876_),
    .A2(_13867_),
    .B1(_13875_),
    .X(_06941_));
 sky130_fd_sc_hd__nand2_1 _18487_ (.A(_13885_),
    .B(_06941_),
    .Y(_06942_));
 sky130_fd_sc_hd__nand4b_1 _18488_ (.A_N(_06919_),
    .B(_13885_),
    .C(_13876_),
    .D(_13868_),
    .Y(_06943_));
 sky130_fd_sc_hd__nor3_1 _18489_ (.A(_13884_),
    .B(_13894_),
    .C(_13903_),
    .Y(_06944_));
 sky130_fd_sc_hd__nand3_1 _18490_ (.A(_06942_),
    .B(_06943_),
    .C(_06944_),
    .Y(_06945_));
 sky130_fd_sc_hd__and2_4 _18491_ (.A(_06940_),
    .B(_06945_),
    .X(_06946_));
 sky130_fd_sc_hd__xor2_2 _18492_ (.A(_13912_),
    .B(_06946_),
    .X(_12534_));
 sky130_fd_sc_hd__inv_1 _18493_ (.A(_12534_),
    .Y(_12700_));
 sky130_fd_sc_hd__clkinv_2 _18494_ (.A(_13908_),
    .Y(_06947_));
 sky130_fd_sc_hd__nor2_1 _18495_ (.A(_13899_),
    .B(_13898_),
    .Y(_06948_));
 sky130_fd_sc_hd__nor2_1 _18496_ (.A(_06947_),
    .B(_06948_),
    .Y(_06949_));
 sky130_fd_sc_hd__nor2_2 _18497_ (.A(_13907_),
    .B(_06949_),
    .Y(_06950_));
 sky130_fd_sc_hd__or3_4 _18498_ (.A(_13888_),
    .B(_13898_),
    .C(_13907_),
    .X(_06951_));
 sky130_fd_sc_hd__a311oi_4 _18499_ (.A1(_13880_),
    .A2(_13889_),
    .A3(_06924_),
    .B1(_06933_),
    .C1(_06951_),
    .Y(_06952_));
 sky130_fd_sc_hd__or2_4 _18500_ (.A(_06950_),
    .B(_06952_),
    .X(_06953_));
 sky130_fd_sc_hd__xnor2_2 _18501_ (.A(_13916_),
    .B(_06953_),
    .Y(_12533_));
 sky130_fd_sc_hd__inv_1 _18502_ (.A(_12533_),
    .Y(_12705_));
 sky130_fd_sc_hd__inv_2 _18503_ (.A(_13920_),
    .Y(_06954_));
 sky130_fd_sc_hd__clkinv_1 _18504_ (.A(_13904_),
    .Y(_06955_));
 sky130_fd_sc_hd__o21bai_4 _18505_ (.A1(_06955_),
    .A2(_06936_),
    .B1_N(_13903_),
    .Y(_06956_));
 sky130_fd_sc_hd__a21oi_2 _18506_ (.A1(_13912_),
    .A2(_06956_),
    .B1(_13911_),
    .Y(_06957_));
 sky130_fd_sc_hd__xnor2_2 _18507_ (.A(_06954_),
    .B(_06957_),
    .Y(_12539_));
 sky130_fd_sc_hd__o21bai_4 _18508_ (.A1(_06938_),
    .A2(_06947_),
    .B1_N(_13907_),
    .Y(_06958_));
 sky130_fd_sc_hd__a21oi_4 _18509_ (.A1(_06958_),
    .A2(_13916_),
    .B1(_13915_),
    .Y(_06959_));
 sky130_fd_sc_hd__xor2_2 _18510_ (.A(_13924_),
    .B(_06959_),
    .X(_12538_));
 sky130_fd_sc_hd__a21oi_1 _18511_ (.A1(_13912_),
    .A2(_06946_),
    .B1(_13911_),
    .Y(_06960_));
 sky130_fd_sc_hd__o21bai_2 _18512_ (.A1(_06954_),
    .A2(_06960_),
    .B1_N(_13919_),
    .Y(_06961_));
 sky130_fd_sc_hd__xor2_2 _18513_ (.A(_13929_),
    .B(_06961_),
    .X(_12544_));
 sky130_fd_sc_hd__clkinv_1 _18514_ (.A(_12544_),
    .Y(_12713_));
 sky130_fd_sc_hd__nor2_1 _18515_ (.A(_06954_),
    .B(_06957_),
    .Y(_06962_));
 sky130_fd_sc_hd__o21ai_0 _18516_ (.A1(_13919_),
    .A2(_06962_),
    .B1(_13929_),
    .Y(_06963_));
 sky130_fd_sc_hd__nand2b_2 _18517_ (.A_N(_13928_),
    .B(_06963_),
    .Y(_06964_));
 sky130_fd_sc_hd__xnor2_2 _18518_ (.A(_13938_),
    .B(_06964_),
    .Y(_12549_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1130 ();
 sky130_fd_sc_hd__nand2_1 _18520_ (.A(_13924_),
    .B(_13933_),
    .Y(_06966_));
 sky130_fd_sc_hd__a21oi_1 _18521_ (.A1(_13933_),
    .A2(_13923_),
    .B1(_13932_),
    .Y(_06967_));
 sky130_fd_sc_hd__o21ai_2 _18522_ (.A1(_06966_),
    .A2(_06959_),
    .B1(_06967_),
    .Y(_06968_));
 sky130_fd_sc_hd__xor2_1 _18523_ (.A(_06968_),
    .B(_13942_),
    .X(_12728_));
 sky130_fd_sc_hd__inv_1 _18524_ (.A(_12728_),
    .Y(_12548_));
 sky130_fd_sc_hd__inv_4 _18525_ (.A(_13947_),
    .Y(_06969_));
 sky130_fd_sc_hd__nand4_1 _18526_ (.A(_13912_),
    .B(_13920_),
    .C(_13929_),
    .D(_13938_),
    .Y(_06970_));
 sky130_fd_sc_hd__inv_1 _18527_ (.A(_06970_),
    .Y(_06971_));
 sky130_fd_sc_hd__a21o_1 _18528_ (.A1(_13920_),
    .A2(_13911_),
    .B1(_13919_),
    .X(_06972_));
 sky130_fd_sc_hd__a21o_1 _18529_ (.A1(_13929_),
    .A2(_06972_),
    .B1(_13928_),
    .X(_06973_));
 sky130_fd_sc_hd__a21o_4 _18530_ (.A1(_13938_),
    .A2(_06973_),
    .B1(_13937_),
    .X(_06974_));
 sky130_fd_sc_hd__a21o_1 _18531_ (.A1(_06946_),
    .A2(_06971_),
    .B1(_06974_),
    .X(_06975_));
 sky130_fd_sc_hd__xnor2_2 _18532_ (.A(_06969_),
    .B(_06975_),
    .Y(_12731_));
 sky130_fd_sc_hd__inv_1 _18533_ (.A(_12731_),
    .Y(_12554_));
 sky130_fd_sc_hd__nor3_2 _18534_ (.A(net345),
    .B(\hash.CA2.e_dash[11] ),
    .C(_06575_),
    .Y(_06976_));
 sky130_fd_sc_hd__a21oi_4 _18535_ (.A1(_06453_),
    .A2(_06575_),
    .B1(_06976_),
    .Y(_13949_));
 sky130_fd_sc_hd__nand4_1 _18536_ (.A(_13924_),
    .B(_13916_),
    .C(_13933_),
    .D(_13942_),
    .Y(_06977_));
 sky130_fd_sc_hd__a21o_1 _18537_ (.A1(_13924_),
    .A2(_13915_),
    .B1(_13923_),
    .X(_06978_));
 sky130_fd_sc_hd__a21o_1 _18538_ (.A1(_13933_),
    .A2(_06978_),
    .B1(_13932_),
    .X(_06979_));
 sky130_fd_sc_hd__a21oi_2 _18539_ (.A1(_13942_),
    .A2(_06979_),
    .B1(_13941_),
    .Y(_06980_));
 sky130_fd_sc_hd__o31ai_4 _18540_ (.A1(_06950_),
    .A2(net1094),
    .A3(_06977_),
    .B1(_06980_),
    .Y(_06981_));
 sky130_fd_sc_hd__xor2_2 _18541_ (.A(_13951_),
    .B(_06981_),
    .X(_12737_));
 sky130_fd_sc_hd__inv_1 _18542_ (.A(_12737_),
    .Y(_12553_));
 sky130_fd_sc_hd__clkinv_2 _18543_ (.A(_13957_),
    .Y(_06982_));
 sky130_fd_sc_hd__nor2_1 _18544_ (.A(_06969_),
    .B(_06982_),
    .Y(_06983_));
 sky130_fd_sc_hd__nor3_1 _18545_ (.A(_06969_),
    .B(_06982_),
    .C(_06970_),
    .Y(_06984_));
 sky130_fd_sc_hd__a222oi_1 _18546_ (.A1(_13957_),
    .A2(_13946_),
    .B1(_06974_),
    .B2(_06983_),
    .C1(_06984_),
    .C2(_06956_),
    .Y(_06985_));
 sky130_fd_sc_hd__nand2b_1 _18547_ (.A_N(_13956_),
    .B(_06985_),
    .Y(_06986_));
 sky130_fd_sc_hd__a21oi_1 _18548_ (.A1(_13966_),
    .A2(_06986_),
    .B1(_13965_),
    .Y(_06987_));
 sky130_fd_sc_hd__xor2_2 _18549_ (.A(_13974_),
    .B(_06987_),
    .X(_12569_));
 sky130_fd_sc_hd__mux2_8 _18550_ (.A0(\hash.CA1.f[14] ),
    .A1(\hash.CA2.e_dash[14] ),
    .S(_06597_),
    .X(_13976_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1129 ();
 sky130_fd_sc_hd__a21o_4 _18552_ (.A1(_13961_),
    .A2(_13950_),
    .B1(_13960_),
    .X(_06989_));
 sky130_fd_sc_hd__inv_1 _18553_ (.A(_13916_),
    .Y(_06990_));
 sky130_fd_sc_hd__nand2_2 _18554_ (.A(_13951_),
    .B(_13961_),
    .Y(_06991_));
 sky130_fd_sc_hd__nand3_1 _18555_ (.A(_13924_),
    .B(_13933_),
    .C(_13942_),
    .Y(_06992_));
 sky130_fd_sc_hd__nor3_1 _18556_ (.A(_06990_),
    .B(_06991_),
    .C(_06992_),
    .Y(_06993_));
 sky130_fd_sc_hd__nor2b_1 _18557_ (.A(_06967_),
    .B_N(_13942_),
    .Y(_06994_));
 sky130_fd_sc_hd__nor2_1 _18558_ (.A(_13941_),
    .B(_06994_),
    .Y(_06995_));
 sky130_fd_sc_hd__nand3_1 _18559_ (.A(_13951_),
    .B(_13961_),
    .C(_13915_),
    .Y(_06996_));
 sky130_fd_sc_hd__o22ai_1 _18560_ (.A1(_06991_),
    .A2(_06995_),
    .B1(_06992_),
    .B2(_06996_),
    .Y(_06997_));
 sky130_fd_sc_hd__a21oi_2 _18561_ (.A1(_06993_),
    .A2(_06958_),
    .B1(_06997_),
    .Y(_06998_));
 sky130_fd_sc_hd__nand2b_1 _18562_ (.A_N(_06989_),
    .B(_06998_),
    .Y(_06999_));
 sky130_fd_sc_hd__a21oi_2 _18563_ (.A1(_06999_),
    .A2(_13970_),
    .B1(_13969_),
    .Y(_07000_));
 sky130_fd_sc_hd__xnor2_2 _18564_ (.A(_07000_),
    .B(_13978_),
    .Y(_12756_));
 sky130_fd_sc_hd__inv_2 _18565_ (.A(_12756_),
    .Y(_12568_));
 sky130_fd_sc_hd__a311o_1 _18566_ (.A1(_06940_),
    .A2(_06945_),
    .A3(_06971_),
    .B1(_06974_),
    .C1(_13946_),
    .X(_07001_));
 sky130_fd_sc_hd__inv_1 _18567_ (.A(_13946_),
    .Y(_07002_));
 sky130_fd_sc_hd__a21oi_2 _18568_ (.A1(_06969_),
    .A2(_07002_),
    .B1(_06982_),
    .Y(_07003_));
 sky130_fd_sc_hd__nor3_2 _18569_ (.A(_13956_),
    .B(_13965_),
    .C(_13973_),
    .Y(_07004_));
 sky130_fd_sc_hd__a21boi_4 _18570_ (.A1(_07001_),
    .A2(_07003_),
    .B1_N(_07004_),
    .Y(_07005_));
 sky130_fd_sc_hd__or2_4 _18571_ (.A(_13966_),
    .B(_13965_),
    .X(_07006_));
 sky130_fd_sc_hd__a21oi_4 _18572_ (.A1(_13974_),
    .A2(_07006_),
    .B1(_13973_),
    .Y(_07007_));
 sky130_fd_sc_hd__nor2_2 _18573_ (.A(_07005_),
    .B(_07007_),
    .Y(_07008_));
 sky130_fd_sc_hd__xnor2_1 _18574_ (.A(_13983_),
    .B(_07008_),
    .Y(_12574_));
 sky130_fd_sc_hd__o21a_1 _18575_ (.A1(_06977_),
    .A2(_06953_),
    .B1(_06980_),
    .X(_07009_));
 sky130_fd_sc_hd__nand3_1 _18576_ (.A(_13951_),
    .B(_13961_),
    .C(_13970_),
    .Y(_07010_));
 sky130_fd_sc_hd__nand2_1 _18577_ (.A(_13970_),
    .B(_06989_),
    .Y(_07011_));
 sky130_fd_sc_hd__o21a_1 _18578_ (.A1(_07010_),
    .A2(_07009_),
    .B1(_07011_),
    .X(_07012_));
 sky130_fd_sc_hd__nand2b_1 _18579_ (.A_N(_13969_),
    .B(_07012_),
    .Y(_07013_));
 sky130_fd_sc_hd__a21oi_2 _18580_ (.A1(_07013_),
    .A2(_13978_),
    .B1(_13977_),
    .Y(_07014_));
 sky130_fd_sc_hd__xnor2_2 _18581_ (.A(_13987_),
    .B(_07014_),
    .Y(_12764_));
 sky130_fd_sc_hd__inv_1 _18582_ (.A(_12764_),
    .Y(_12573_));
 sky130_fd_sc_hd__nor3_1 _18583_ (.A(net342),
    .B(\hash.CA2.e_dash[16] ),
    .C(\hash.CA1.S1.X[16] ),
    .Y(_07015_));
 sky130_fd_sc_hd__a21oi_4 _18584_ (.A1(_06462_),
    .A2(\hash.CA1.S1.X[16] ),
    .B1(_07015_),
    .Y(_13995_));
 sky130_fd_sc_hd__inv_6 _18585_ (.A(_06568_),
    .Y(\hash.CA1.S1.X[10] ));
 sky130_fd_sc_hd__mux2_8 _18586_ (.A0(_06467_),
    .A1(\hash.CA2.e_dash[18] ),
    .S(_06634_),
    .X(_14012_));
 sky130_fd_sc_hd__and4_4 _18587_ (.A(_13983_),
    .B(_13993_),
    .C(_14002_),
    .D(_14010_),
    .X(_07016_));
 sky130_fd_sc_hd__nand3_1 _18588_ (.A(_14018_),
    .B(_14026_),
    .C(_07016_),
    .Y(_07017_));
 sky130_fd_sc_hd__a211oi_2 _18589_ (.A1(_06985_),
    .A2(_07004_),
    .B1(_07007_),
    .C1(_07017_),
    .Y(_07018_));
 sky130_fd_sc_hd__a21o_1 _18590_ (.A1(_13993_),
    .A2(_13982_),
    .B1(_13992_),
    .X(_07019_));
 sky130_fd_sc_hd__a21o_1 _18591_ (.A1(_14002_),
    .A2(_07019_),
    .B1(_14001_),
    .X(_07020_));
 sky130_fd_sc_hd__a21o_4 _18592_ (.A1(_14010_),
    .A2(_07020_),
    .B1(_14009_),
    .X(_07021_));
 sky130_fd_sc_hd__a21oi_1 _18593_ (.A1(_14018_),
    .A2(_07021_),
    .B1(_14017_),
    .Y(_07022_));
 sky130_fd_sc_hd__nor2b_2 _18594_ (.A(_07022_),
    .B_N(_14026_),
    .Y(_07023_));
 sky130_fd_sc_hd__a21oi_2 _18595_ (.A1(_06985_),
    .A2(_07004_),
    .B1(_07007_),
    .Y(_07024_));
 sky130_fd_sc_hd__and2_0 _18596_ (.A(_07024_),
    .B(_07016_),
    .X(_07025_));
 sky130_fd_sc_hd__o21ai_0 _18597_ (.A1(_07025_),
    .A2(_07021_),
    .B1(_14018_),
    .Y(_07026_));
 sky130_fd_sc_hd__nor3b_1 _18598_ (.A(_14026_),
    .B(_14017_),
    .C_N(_07026_),
    .Y(_07027_));
 sky130_fd_sc_hd__nor3_2 _18599_ (.A(_07018_),
    .B(_07023_),
    .C(_07027_),
    .Y(_12599_));
 sky130_fd_sc_hd__clkinv_2 _18600_ (.A(_12599_),
    .Y(_12792_));
 sky130_fd_sc_hd__a21o_1 _18601_ (.A1(_14026_),
    .A2(_14017_),
    .B1(_14025_),
    .X(_07028_));
 sky130_fd_sc_hd__nand2_1 _18602_ (.A(_14018_),
    .B(_14026_),
    .Y(_07029_));
 sky130_fd_sc_hd__a21oi_1 _18603_ (.A1(_07008_),
    .A2(_07016_),
    .B1(_07021_),
    .Y(_07030_));
 sky130_fd_sc_hd__nor2_1 _18604_ (.A(_07029_),
    .B(_07030_),
    .Y(_07031_));
 sky130_fd_sc_hd__nor2_1 _18605_ (.A(_07028_),
    .B(_07031_),
    .Y(_07032_));
 sky130_fd_sc_hd__xnor2_1 _18606_ (.A(_14034_),
    .B(_07032_),
    .Y(_12801_));
 sky130_fd_sc_hd__inv_1 _18607_ (.A(_12801_),
    .Y(_12604_));
 sky130_fd_sc_hd__nand2_4 _18608_ (.A(_13997_),
    .B(_14006_),
    .Y(_07033_));
 sky130_fd_sc_hd__nand2_1 _18609_ (.A(_13978_),
    .B(_13987_),
    .Y(_07034_));
 sky130_fd_sc_hd__nor2_1 _18610_ (.A(_07010_),
    .B(_07034_),
    .Y(_07035_));
 sky130_fd_sc_hd__a21o_1 _18611_ (.A1(_13978_),
    .A2(_13969_),
    .B1(_13977_),
    .X(_07036_));
 sky130_fd_sc_hd__a21oi_1 _18612_ (.A1(_13987_),
    .A2(_07036_),
    .B1(_13986_),
    .Y(_07037_));
 sky130_fd_sc_hd__o21ai_0 _18613_ (.A1(_07011_),
    .A2(_07034_),
    .B1(_07037_),
    .Y(_07038_));
 sky130_fd_sc_hd__a21oi_2 _18614_ (.A1(_06981_),
    .A2(_07035_),
    .B1(_07038_),
    .Y(_07039_));
 sky130_fd_sc_hd__nand2_4 _18615_ (.A(_14006_),
    .B(_13996_),
    .Y(_07040_));
 sky130_fd_sc_hd__o21ai_4 _18616_ (.A1(_07033_),
    .A2(_07039_),
    .B1(_07040_),
    .Y(_07041_));
 sky130_fd_sc_hd__and3_4 _18617_ (.A(_14014_),
    .B(_14022_),
    .C(_14030_),
    .X(_07042_));
 sky130_fd_sc_hd__a21o_1 _18618_ (.A1(_14014_),
    .A2(_14005_),
    .B1(_14013_),
    .X(_07043_));
 sky130_fd_sc_hd__a21o_1 _18619_ (.A1(_14022_),
    .A2(_07043_),
    .B1(_14021_),
    .X(_07044_));
 sky130_fd_sc_hd__a21o_1 _18620_ (.A1(_14030_),
    .A2(_07044_),
    .B1(_14029_),
    .X(_07045_));
 sky130_fd_sc_hd__a21o_1 _18621_ (.A1(_07041_),
    .A2(_07042_),
    .B1(_07045_),
    .X(_07046_));
 sky130_fd_sc_hd__xor2_1 _18622_ (.A(_14038_),
    .B(_07046_),
    .X(_12807_));
 sky130_fd_sc_hd__inv_1 _18623_ (.A(_12807_),
    .Y(_12603_));
 sky130_fd_sc_hd__o31ai_1 _18624_ (.A1(_14025_),
    .A2(_07018_),
    .A3(_07023_),
    .B1(_14034_),
    .Y(_07047_));
 sky130_fd_sc_hd__nor2_1 _18625_ (.A(_14043_),
    .B(_14033_),
    .Y(_07048_));
 sky130_fd_sc_hd__o21a_1 _18626_ (.A1(_14034_),
    .A2(_14033_),
    .B1(_14043_),
    .X(_07049_));
 sky130_fd_sc_hd__o41a_1 _18627_ (.A1(_14025_),
    .A2(_14033_),
    .A3(_07018_),
    .A4(_07023_),
    .B1(_07049_),
    .X(_07050_));
 sky130_fd_sc_hd__a21o_4 _18628_ (.A1(_07047_),
    .A2(_07048_),
    .B1(_07050_),
    .X(_12609_));
 sky130_fd_sc_hd__nor3_1 _18629_ (.A(_13969_),
    .B(_13977_),
    .C(_06989_),
    .Y(_07051_));
 sky130_fd_sc_hd__or2_0 _18630_ (.A(_13970_),
    .B(_13969_),
    .X(_07052_));
 sky130_fd_sc_hd__a21oi_1 _18631_ (.A1(_13978_),
    .A2(_07052_),
    .B1(_13977_),
    .Y(_07053_));
 sky130_fd_sc_hd__a21oi_2 _18632_ (.A1(_07051_),
    .A2(_06998_),
    .B1(_07053_),
    .Y(_07054_));
 sky130_fd_sc_hd__a21oi_4 _18633_ (.A1(_07054_),
    .A2(_13987_),
    .B1(_13986_),
    .Y(_07055_));
 sky130_fd_sc_hd__o21ai_4 _18634_ (.A1(_07055_),
    .A2(_07033_),
    .B1(_07040_),
    .Y(_07056_));
 sky130_fd_sc_hd__a21o_1 _18635_ (.A1(_14038_),
    .A2(_07045_),
    .B1(_14037_),
    .X(_07057_));
 sky130_fd_sc_hd__a31o_1 _18636_ (.A1(_14038_),
    .A2(_07042_),
    .A3(_07056_),
    .B1(_07057_),
    .X(_07058_));
 sky130_fd_sc_hd__xor2_1 _18637_ (.A(_14047_),
    .B(_07058_),
    .X(_12814_));
 sky130_fd_sc_hd__inv_1 _18638_ (.A(_12814_),
    .Y(_12608_));
 sky130_fd_sc_hd__and3_1 _18639_ (.A(_14018_),
    .B(_14026_),
    .C(_14034_),
    .X(_07059_));
 sky130_fd_sc_hd__nand3_1 _18640_ (.A(_14043_),
    .B(_07016_),
    .C(_07059_),
    .Y(_07060_));
 sky130_fd_sc_hd__nand2_1 _18641_ (.A(_07021_),
    .B(_07059_),
    .Y(_07061_));
 sky130_fd_sc_hd__a21oi_1 _18642_ (.A1(_14034_),
    .A2(_07028_),
    .B1(_14033_),
    .Y(_07062_));
 sky130_fd_sc_hd__a21bo_1 _18643_ (.A1(_07061_),
    .A2(_07062_),
    .B1_N(_14043_),
    .X(_07063_));
 sky130_fd_sc_hd__clkinv_1 _18644_ (.A(_14042_),
    .Y(_07064_));
 sky130_fd_sc_hd__o311ai_2 _18645_ (.A1(_07005_),
    .A2(_07007_),
    .A3(_07060_),
    .B1(_07063_),
    .C1(_07064_),
    .Y(_07065_));
 sky130_fd_sc_hd__xor2_2 _18646_ (.A(_14053_),
    .B(_07065_),
    .X(_12817_));
 sky130_fd_sc_hd__inv_1 _18647_ (.A(_12817_),
    .Y(_12614_));
 sky130_fd_sc_hd__nand3_2 _18648_ (.A(_14038_),
    .B(_14047_),
    .C(_07042_),
    .Y(_07066_));
 sky130_fd_sc_hd__nor2b_1 _18649_ (.A(_07066_),
    .B_N(_07041_),
    .Y(_07067_));
 sky130_fd_sc_hd__a21oi_2 _18650_ (.A1(_14047_),
    .A2(_07057_),
    .B1(_14046_),
    .Y(_07068_));
 sky130_fd_sc_hd__nor2b_1 _18651_ (.A(_07067_),
    .B_N(_07068_),
    .Y(_07069_));
 sky130_fd_sc_hd__xnor2_1 _18652_ (.A(_14057_),
    .B(_07069_),
    .Y(_12823_));
 sky130_fd_sc_hd__inv_1 _18653_ (.A(_12823_),
    .Y(_12613_));
 sky130_fd_sc_hd__o21ai_0 _18654_ (.A1(_14042_),
    .A2(_07050_),
    .B1(_14053_),
    .Y(_07070_));
 sky130_fd_sc_hd__nand2b_2 _18655_ (.A_N(_14052_),
    .B(_07070_),
    .Y(_07071_));
 sky130_fd_sc_hd__xnor2_2 _18656_ (.A(_14063_),
    .B(_07071_),
    .Y(_12619_));
 sky130_fd_sc_hd__mux2_1 _18657_ (.A0(_06487_),
    .A1(\hash.CA2.e_dash[24] ),
    .S(_06673_),
    .X(_14065_));
 sky130_fd_sc_hd__inv_1 _18658_ (.A(_07056_),
    .Y(_07072_));
 sky130_fd_sc_hd__o21ai_0 _18659_ (.A1(_07072_),
    .A2(_07066_),
    .B1(_07068_),
    .Y(_07073_));
 sky130_fd_sc_hd__a21oi_1 _18660_ (.A1(_14057_),
    .A2(_07073_),
    .B1(_14056_),
    .Y(_07074_));
 sky130_fd_sc_hd__xnor2_1 _18661_ (.A(_07074_),
    .B(_14067_),
    .Y(_12830_));
 sky130_fd_sc_hd__inv_1 _18662_ (.A(_12830_),
    .Y(_12618_));
 sky130_fd_sc_hd__a21o_1 _18663_ (.A1(_14053_),
    .A2(_07065_),
    .B1(_14052_),
    .X(_07075_));
 sky130_fd_sc_hd__a21o_4 _18664_ (.A1(_14063_),
    .A2(_07075_),
    .B1(_14062_),
    .X(_07076_));
 sky130_fd_sc_hd__xor2_2 _18665_ (.A(_14073_),
    .B(_07076_),
    .X(_12833_));
 sky130_fd_sc_hd__inv_1 _18666_ (.A(_12833_),
    .Y(_12624_));
 sky130_fd_sc_hd__nor3_1 _18667_ (.A(net534),
    .B(\hash.CA2.e_dash[25] ),
    .C(_06683_),
    .Y(_07077_));
 sky130_fd_sc_hd__a21oi_4 _18668_ (.A1(_06490_),
    .A2(_06683_),
    .B1(_07077_),
    .Y(_14075_));
 sky130_fd_sc_hd__clkinv_1 _18669_ (.A(_14077_),
    .Y(_07078_));
 sky130_fd_sc_hd__nand2_2 _18670_ (.A(_14067_),
    .B(_14057_),
    .Y(_07079_));
 sky130_fd_sc_hd__nor2_2 _18671_ (.A(_07066_),
    .B(_07079_),
    .Y(_07080_));
 sky130_fd_sc_hd__nand2_1 _18672_ (.A(_14067_),
    .B(_14056_),
    .Y(_07081_));
 sky130_fd_sc_hd__o21ai_2 _18673_ (.A1(_07068_),
    .A2(_07079_),
    .B1(_07081_),
    .Y(_07082_));
 sky130_fd_sc_hd__a211o_4 _18674_ (.A1(_07041_),
    .A2(_07080_),
    .B1(_07082_),
    .C1(_14066_),
    .X(_07083_));
 sky130_fd_sc_hd__xnor2_1 _18675_ (.A(_07078_),
    .B(_07083_),
    .Y(_12839_));
 sky130_fd_sc_hd__inv_1 _18676_ (.A(_12839_),
    .Y(_12623_));
 sky130_fd_sc_hd__nand2_1 _18677_ (.A(_14073_),
    .B(_07076_),
    .Y(_07084_));
 sky130_fd_sc_hd__nand2b_1 _18678_ (.A_N(_14072_),
    .B(_07084_),
    .Y(_07085_));
 sky130_fd_sc_hd__a21o_1 _18679_ (.A1(_14083_),
    .A2(_07085_),
    .B1(_14082_),
    .X(_07086_));
 sky130_fd_sc_hd__xor2_2 _18680_ (.A(_14092_),
    .B(_07086_),
    .X(_12848_));
 sky130_fd_sc_hd__inv_1 _18681_ (.A(_12848_),
    .Y(_12634_));
 sky130_fd_sc_hd__nor3_1 _18682_ (.A(net534),
    .B(\hash.CA2.e_dash[27] ),
    .C(net1124),
    .Y(_07087_));
 sky130_fd_sc_hd__a21oi_2 _18683_ (.A1(_06497_),
    .A2(net1124),
    .B1(_07087_),
    .Y(_14094_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1128 ();
 sky130_fd_sc_hd__a21o_1 _18685_ (.A1(_14077_),
    .A2(_07083_),
    .B1(_14076_),
    .X(_07089_));
 sky130_fd_sc_hd__a21oi_1 _18686_ (.A1(_14087_),
    .A2(_07089_),
    .B1(_14086_),
    .Y(_07090_));
 sky130_fd_sc_hd__xnor2_1 _18687_ (.A(_14096_),
    .B(_07090_),
    .Y(_12853_));
 sky130_fd_sc_hd__inv_1 _18688_ (.A(_12853_),
    .Y(_12633_));
 sky130_fd_sc_hd__o211ai_1 _18689_ (.A1(_14042_),
    .A2(_07050_),
    .B1(_14053_),
    .C1(_14063_),
    .Y(_07091_));
 sky130_fd_sc_hd__a21oi_1 _18690_ (.A1(_14063_),
    .A2(_14052_),
    .B1(_14062_),
    .Y(_07092_));
 sky130_fd_sc_hd__a21boi_2 _18691_ (.A1(_07091_),
    .A2(_07092_),
    .B1_N(_14073_),
    .Y(_07093_));
 sky130_fd_sc_hd__o21ai_0 _18692_ (.A1(_14083_),
    .A2(_14082_),
    .B1(_14092_),
    .Y(_07094_));
 sky130_fd_sc_hd__nand2b_1 _18693_ (.A_N(_14091_),
    .B(_07094_),
    .Y(_07095_));
 sky130_fd_sc_hd__o41ai_2 _18694_ (.A1(_14072_),
    .A2(_14082_),
    .A3(_14091_),
    .A4(_07093_),
    .B1(_07095_),
    .Y(_07096_));
 sky130_fd_sc_hd__xnor2_2 _18695_ (.A(_14101_),
    .B(_07096_),
    .Y(_12856_));
 sky130_fd_sc_hd__inv_1 _18696_ (.A(_12856_),
    .Y(_12639_));
 sky130_fd_sc_hd__nor2_1 _18697_ (.A(\hash.CA2.e_dash[28] ),
    .B(_06707_),
    .Y(_07097_));
 sky130_fd_sc_hd__a31oi_2 _18698_ (.A1(_06002_),
    .A2(_06501_),
    .A3(_06707_),
    .B1(_07097_),
    .Y(_14103_));
 sky130_fd_sc_hd__a211oi_4 _18699_ (.A1(_07056_),
    .A2(_07080_),
    .B1(_07082_),
    .C1(_14066_),
    .Y(_07098_));
 sky130_fd_sc_hd__nand2_1 _18700_ (.A(_14077_),
    .B(_14087_),
    .Y(_07099_));
 sky130_fd_sc_hd__a21oi_1 _18701_ (.A1(_14087_),
    .A2(_14076_),
    .B1(_14086_),
    .Y(_07100_));
 sky130_fd_sc_hd__o21ai_1 _18702_ (.A1(_07098_),
    .A2(_07099_),
    .B1(_07100_),
    .Y(_07101_));
 sky130_fd_sc_hd__a21o_1 _18703_ (.A1(_14096_),
    .A2(_07101_),
    .B1(_14095_),
    .X(_07102_));
 sky130_fd_sc_hd__xor2_2 _18704_ (.A(_14105_),
    .B(_07102_),
    .X(_12861_));
 sky130_fd_sc_hd__inv_1 _18705_ (.A(_12861_),
    .Y(_12638_));
 sky130_fd_sc_hd__nand2_1 _18706_ (.A(_14101_),
    .B(_14111_),
    .Y(_07103_));
 sky130_fd_sc_hd__inv_1 _18707_ (.A(_14101_),
    .Y(_07104_));
 sky130_fd_sc_hd__nor3b_1 _18708_ (.A(_14100_),
    .B(_14110_),
    .C_N(_14120_),
    .Y(_07105_));
 sky130_fd_sc_hd__o21ai_0 _18709_ (.A1(_07104_),
    .A2(_07096_),
    .B1(_07105_),
    .Y(_07106_));
 sky130_fd_sc_hd__o31ai_1 _18710_ (.A1(_14120_),
    .A2(_07096_),
    .A3(_07103_),
    .B1(_07106_),
    .Y(_07107_));
 sky130_fd_sc_hd__a21oi_1 _18711_ (.A1(_14111_),
    .A2(_14100_),
    .B1(_14110_),
    .Y(_07108_));
 sky130_fd_sc_hd__nor2_1 _18712_ (.A(_14120_),
    .B(_07108_),
    .Y(_07109_));
 sky130_fd_sc_hd__nor3b_1 _18713_ (.A(_14111_),
    .B(_14110_),
    .C_N(_14120_),
    .Y(_07110_));
 sky130_fd_sc_hd__nor3_2 _18714_ (.A(_07107_),
    .B(_07109_),
    .C(_07110_),
    .Y(_12649_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1127 ();
 sky130_fd_sc_hd__nand4_1 _18716_ (.A(_14096_),
    .B(_14105_),
    .C(_14115_),
    .D(_07101_),
    .Y(_07112_));
 sky130_fd_sc_hd__nand2_1 _18717_ (.A(_14115_),
    .B(_14104_),
    .Y(_07113_));
 sky130_fd_sc_hd__nand3_1 _18718_ (.A(_14105_),
    .B(_14115_),
    .C(_14095_),
    .Y(_07114_));
 sky130_fd_sc_hd__nand4b_1 _18719_ (.A_N(_14114_),
    .B(_07112_),
    .C(_07113_),
    .D(_07114_),
    .Y(_07115_));
 sky130_fd_sc_hd__xnor2_1 _18720_ (.A(_14124_),
    .B(_07115_),
    .Y(_12648_));
 sky130_fd_sc_hd__o21bai_4 _18721_ (.A1(_06990_),
    .A2(_06953_),
    .B1_N(_13915_),
    .Y(_07116_));
 sky130_fd_sc_hd__a21oi_4 _18722_ (.A1(_13924_),
    .A2(_07116_),
    .B1(_13923_),
    .Y(_07117_));
 sky130_fd_sc_hd__xnor2_2 _18723_ (.A(_13933_),
    .B(_07117_),
    .Y(_12720_));
 sky130_fd_sc_hd__o21ai_1 _18724_ (.A1(_06959_),
    .A2(_06992_),
    .B1(_06995_),
    .Y(_07118_));
 sky130_fd_sc_hd__a21oi_2 _18725_ (.A1(_07118_),
    .A2(_13951_),
    .B1(_13950_),
    .Y(_07119_));
 sky130_fd_sc_hd__xnor2_1 _18726_ (.A(_13961_),
    .B(_07119_),
    .Y(_12743_));
 sky130_fd_sc_hd__nor2_1 _18727_ (.A(_07009_),
    .B(_06991_),
    .Y(_07120_));
 sky130_fd_sc_hd__o31a_1 _18728_ (.A1(_13970_),
    .A2(_06989_),
    .A3(_07120_),
    .B1(_07012_),
    .X(_12749_));
 sky130_fd_sc_hd__xnor2_1 _18729_ (.A(_13997_),
    .B(_07055_),
    .Y(_12771_));
 sky130_fd_sc_hd__nor2_1 _18730_ (.A(_14006_),
    .B(_13996_),
    .Y(_07121_));
 sky130_fd_sc_hd__nand2b_1 _18731_ (.A_N(_07039_),
    .B(_13997_),
    .Y(_07122_));
 sky130_fd_sc_hd__a21oi_1 _18732_ (.A1(_07121_),
    .A2(_07122_),
    .B1(_07041_),
    .Y(_12777_));
 sky130_fd_sc_hd__nor2_2 _18733_ (.A(_14005_),
    .B(_07056_),
    .Y(_07123_));
 sky130_fd_sc_hd__xnor2_1 _18734_ (.A(_14014_),
    .B(_07123_),
    .Y(_12783_));
 sky130_fd_sc_hd__o21a_1 _18735_ (.A1(_14005_),
    .A2(_07041_),
    .B1(_14014_),
    .X(_07124_));
 sky130_fd_sc_hd__nor2_2 _18736_ (.A(_14013_),
    .B(_07124_),
    .Y(_07125_));
 sky130_fd_sc_hd__xnor2_1 _18737_ (.A(_14022_),
    .B(_07125_),
    .Y(_12789_));
 sky130_fd_sc_hd__o21ai_0 _18738_ (.A1(_14005_),
    .A2(_07056_),
    .B1(_14014_),
    .Y(_07126_));
 sky130_fd_sc_hd__nand2b_1 _18739_ (.A_N(_14013_),
    .B(_07126_),
    .Y(_07127_));
 sky130_fd_sc_hd__a21oi_2 _18740_ (.A1(_14022_),
    .A2(_07127_),
    .B1(_14021_),
    .Y(_07128_));
 sky130_fd_sc_hd__xnor2_1 _18741_ (.A(_14030_),
    .B(_07128_),
    .Y(_12798_));
 sky130_fd_sc_hd__o21bai_2 _18742_ (.A1(_07078_),
    .A2(_07098_),
    .B1_N(_14076_),
    .Y(_07129_));
 sky130_fd_sc_hd__xor2_1 _18743_ (.A(_14087_),
    .B(_07129_),
    .X(_12845_));
 sky130_fd_sc_hd__a2111o_1 _18744_ (.A1(_14077_),
    .A2(_07083_),
    .B1(_14095_),
    .C1(_14086_),
    .D1(_14076_),
    .X(_07130_));
 sky130_fd_sc_hd__nor3_1 _18745_ (.A(_14087_),
    .B(_14086_),
    .C(_14095_),
    .Y(_07131_));
 sky130_fd_sc_hd__nor2_1 _18746_ (.A(_14096_),
    .B(_14095_),
    .Y(_07132_));
 sky130_fd_sc_hd__nor2_1 _18747_ (.A(_07131_),
    .B(_07132_),
    .Y(_07133_));
 sky130_fd_sc_hd__a31oi_2 _18748_ (.A1(_14105_),
    .A2(_07130_),
    .A3(_07133_),
    .B1(_14104_),
    .Y(_07134_));
 sky130_fd_sc_hd__xnor2_1 _18749_ (.A(_14115_),
    .B(_07134_),
    .Y(_12867_));
 sky130_fd_sc_hd__clkinvlp_4 _18750_ (.A(net1037),
    .Y(_00906_));
 sky130_fd_sc_hd__inv_1 _18751_ (.A(_12988_),
    .Y(_11600_));
 sky130_fd_sc_hd__inv_1 _18752_ (.A(_13111_),
    .Y(_11848_));
 sky130_fd_sc_hd__clkinv_2 _18753_ (.A(_13231_),
    .Y(_12083_));
 sky130_fd_sc_hd__inv_1 _18754_ (.A(_13240_),
    .Y(_12105_));
 sky130_fd_sc_hd__inv_1 _18755_ (.A(\hash.CA1.k_i2[1] ),
    .Y(_12366_));
 sky130_fd_sc_hd__inv_2 _18756_ (.A(\hash.CA1.k_i2[0] ),
    .Y(_12371_));
 sky130_fd_sc_hd__clkinv_1 _18757_ (.A(\hash.CA1.k_i2[3] ),
    .Y(_12381_));
 sky130_fd_sc_hd__clkinv_1 _18758_ (.A(\hash.CA1.k_i2[5] ),
    .Y(_12389_));
 sky130_fd_sc_hd__inv_1 _18759_ (.A(\hash.CA1.k_i2[7] ),
    .Y(_12397_));
 sky130_fd_sc_hd__inv_2 _18760_ (.A(\hash.CA1.k_i2[8] ),
    .Y(_12402_));
 sky130_fd_sc_hd__inv_2 _18761_ (.A(\hash.CA1.k_i2[11] ),
    .Y(_12413_));
 sky130_fd_sc_hd__inv_2 _18762_ (.A(\hash.CA1.k_i2[12] ),
    .Y(_12418_));
 sky130_fd_sc_hd__inv_1 _18763_ (.A(\hash.CA1.k_i2[14] ),
    .Y(_12426_));
 sky130_fd_sc_hd__inv_1 _18764_ (.A(\hash.CA1.k_i2[15] ),
    .Y(_12431_));
 sky130_fd_sc_hd__inv_1 _18765_ (.A(\hash.CA1.k_i2[16] ),
    .Y(_12436_));
 sky130_fd_sc_hd__inv_1 _18766_ (.A(\hash.CA1.k_i2[17] ),
    .Y(_12441_));
 sky130_fd_sc_hd__inv_2 _18767_ (.A(\hash.CA1.k_i2[23] ),
    .Y(_12461_));
 sky130_fd_sc_hd__inv_2 _18768_ (.A(\hash.CA1.k_i2[24] ),
    .Y(_12466_));
 sky130_fd_sc_hd__inv_1 _18769_ (.A(\hash.CA1.k_i2[25] ),
    .Y(_12471_));
 sky130_fd_sc_hd__inv_1 _18770_ (.A(\hash.CA1.k_i2[26] ),
    .Y(_12476_));
 sky130_fd_sc_hd__inv_1 _18771_ (.A(\hash.CA1.k_i2[27] ),
    .Y(_12481_));
 sky130_fd_sc_hd__inv_1 _18772_ (.A(\hash.CA1.k_i2[28] ),
    .Y(_12486_));
 sky130_fd_sc_hd__clkinv_1 _18773_ (.A(_12724_),
    .Y(_12736_));
 sky130_fd_sc_hd__inv_1 _18774_ (.A(_14204_),
    .Y(_12879_));
 sky130_fd_sc_hd__inv_1 _18775_ (.A(_14207_),
    .Y(_12884_));
 sky130_fd_sc_hd__inv_1 _18776_ (.A(_14208_),
    .Y(_12889_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1123 ();
 sky130_fd_sc_hd__mux4_2 _18781_ (.A0(\w[1][0] ),
    .A1(\w[5][0] ),
    .A2(\w[3][0] ),
    .A3(\w[7][0] ),
    .S0(net401),
    .S1(net408),
    .X(_07139_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1119 ();
 sky130_fd_sc_hd__mux4_2 _18786_ (.A0(\w[9][0] ),
    .A1(\w[13][0] ),
    .A2(\w[11][0] ),
    .A3(\w[15][0] ),
    .S0(net401),
    .S1(net408),
    .X(_07144_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1117 ();
 sky130_fd_sc_hd__mux4_2 _18789_ (.A0(\w[17][0] ),
    .A1(\w[21][0] ),
    .A2(\w[19][0] ),
    .A3(\w[23][0] ),
    .S0(net401),
    .S1(net408),
    .X(_07147_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1114 ();
 sky130_fd_sc_hd__mux4_2 _18793_ (.A0(\w[25][0] ),
    .A1(\w[29][0] ),
    .A2(\w[27][0] ),
    .A3(\w[31][0] ),
    .S0(net401),
    .S1(net408),
    .X(_07151_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1110 ();
 sky130_fd_sc_hd__mux4_2 _18798_ (.A0(_07139_),
    .A1(_07144_),
    .A2(_07147_),
    .A3(_07151_),
    .S0(net398),
    .S1(net396),
    .X(_07156_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1108 ();
 sky130_fd_sc_hd__mux4_2 _18801_ (.A0(\w[33][0] ),
    .A1(\w[37][0] ),
    .A2(\w[35][0] ),
    .A3(\w[39][0] ),
    .S0(net406),
    .S1(net408),
    .X(_07159_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1106 ();
 sky130_fd_sc_hd__mux4_2 _18804_ (.A0(\w[41][0] ),
    .A1(\w[45][0] ),
    .A2(\w[43][0] ),
    .A3(\w[47][0] ),
    .S0(net406),
    .S1(net408),
    .X(_07162_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1104 ();
 sky130_fd_sc_hd__mux4_2 _18807_ (.A0(\w[49][0] ),
    .A1(\w[53][0] ),
    .A2(\w[51][0] ),
    .A3(\w[55][0] ),
    .S0(net406),
    .S1(net408),
    .X(_07165_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1102 ();
 sky130_fd_sc_hd__mux4_2 _18810_ (.A0(\w[57][0] ),
    .A1(\w[61][0] ),
    .A2(\w[59][0] ),
    .A3(\w[63][0] ),
    .S0(net406),
    .S1(net408),
    .X(_07168_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1100 ();
 sky130_fd_sc_hd__mux4_2 _18813_ (.A0(_07159_),
    .A1(_07162_),
    .A2(_07165_),
    .A3(_07168_),
    .S0(net398),
    .S1(net396),
    .X(_07171_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1099 ();
 sky130_fd_sc_hd__mux2i_4 _18815_ (.A0(_07156_),
    .A1(_07171_),
    .S(net394),
    .Y(_11580_));
 sky130_fd_sc_hd__mux4_2 _18816_ (.A0(\w[1][1] ),
    .A1(\w[5][1] ),
    .A2(\w[3][1] ),
    .A3(\w[7][1] ),
    .S0(net401),
    .S1(net408),
    .X(_07173_));
 sky130_fd_sc_hd__mux4_2 _18817_ (.A0(\w[9][1] ),
    .A1(\w[13][1] ),
    .A2(\w[11][1] ),
    .A3(\w[15][1] ),
    .S0(net401),
    .S1(net408),
    .X(_07174_));
 sky130_fd_sc_hd__mux4_2 _18818_ (.A0(\w[17][1] ),
    .A1(\w[21][1] ),
    .A2(\w[19][1] ),
    .A3(\w[23][1] ),
    .S0(net401),
    .S1(net408),
    .X(_07175_));
 sky130_fd_sc_hd__mux4_2 _18819_ (.A0(\w[25][1] ),
    .A1(\w[29][1] ),
    .A2(\w[27][1] ),
    .A3(\w[31][1] ),
    .S0(net401),
    .S1(net408),
    .X(_07176_));
 sky130_fd_sc_hd__mux4_2 _18820_ (.A0(_07173_),
    .A1(_07174_),
    .A2(_07175_),
    .A3(_07176_),
    .S0(net398),
    .S1(net396),
    .X(_07177_));
 sky130_fd_sc_hd__mux4_2 _18821_ (.A0(\w[33][1] ),
    .A1(\w[37][1] ),
    .A2(\w[35][1] ),
    .A3(\w[39][1] ),
    .S0(net401),
    .S1(net408),
    .X(_07178_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1098 ();
 sky130_fd_sc_hd__mux4_2 _18823_ (.A0(\w[41][1] ),
    .A1(\w[45][1] ),
    .A2(\w[43][1] ),
    .A3(\w[47][1] ),
    .S0(net405),
    .S1(net408),
    .X(_07180_));
 sky130_fd_sc_hd__mux4_2 _18824_ (.A0(\w[49][1] ),
    .A1(\w[53][1] ),
    .A2(\w[51][1] ),
    .A3(\w[55][1] ),
    .S0(net401),
    .S1(net408),
    .X(_07181_));
 sky130_fd_sc_hd__mux4_2 _18825_ (.A0(\w[57][1] ),
    .A1(\w[61][1] ),
    .A2(\w[59][1] ),
    .A3(\w[63][1] ),
    .S0(net405),
    .S1(net408),
    .X(_07182_));
 sky130_fd_sc_hd__mux4_2 _18826_ (.A0(_07178_),
    .A1(_07180_),
    .A2(_07181_),
    .A3(_07182_),
    .S0(net398),
    .S1(net536),
    .X(_07183_));
 sky130_fd_sc_hd__mux2i_4 _18827_ (.A0(_07177_),
    .A1(_07183_),
    .S(net395),
    .Y(_11585_));
 sky130_fd_sc_hd__mux4_2 _18828_ (.A0(\w[1][2] ),
    .A1(\w[5][2] ),
    .A2(\w[3][2] ),
    .A3(\w[7][2] ),
    .S0(net401),
    .S1(net408),
    .X(_07184_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1097 ();
 sky130_fd_sc_hd__mux4_2 _18830_ (.A0(\w[9][2] ),
    .A1(\w[13][2] ),
    .A2(\w[11][2] ),
    .A3(\w[15][2] ),
    .S0(net401),
    .S1(net408),
    .X(_07186_));
 sky130_fd_sc_hd__mux4_2 _18831_ (.A0(\w[17][2] ),
    .A1(\w[21][2] ),
    .A2(\w[19][2] ),
    .A3(\w[23][2] ),
    .S0(net401),
    .S1(net408),
    .X(_07187_));
 sky130_fd_sc_hd__mux4_2 _18832_ (.A0(\w[25][2] ),
    .A1(\w[29][2] ),
    .A2(\w[27][2] ),
    .A3(\w[31][2] ),
    .S0(net401),
    .S1(net408),
    .X(_07188_));
 sky130_fd_sc_hd__mux4_2 _18833_ (.A0(_07184_),
    .A1(_07186_),
    .A2(_07187_),
    .A3(_07188_),
    .S0(net398),
    .S1(net396),
    .X(_07189_));
 sky130_fd_sc_hd__mux4_2 _18834_ (.A0(\w[33][2] ),
    .A1(\w[37][2] ),
    .A2(\w[35][2] ),
    .A3(\w[39][2] ),
    .S0(net404),
    .S1(net411),
    .X(_07190_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1096 ();
 sky130_fd_sc_hd__mux4_2 _18836_ (.A0(\w[41][2] ),
    .A1(\w[45][2] ),
    .A2(\w[43][2] ),
    .A3(\w[47][2] ),
    .S0(net404),
    .S1(net411),
    .X(_07192_));
 sky130_fd_sc_hd__mux4_2 _18837_ (.A0(\w[49][2] ),
    .A1(\w[53][2] ),
    .A2(\w[51][2] ),
    .A3(\w[55][2] ),
    .S0(net404),
    .S1(net411),
    .X(_07193_));
 sky130_fd_sc_hd__mux4_2 _18838_ (.A0(\w[57][2] ),
    .A1(\w[61][2] ),
    .A2(\w[59][2] ),
    .A3(\w[63][2] ),
    .S0(net403),
    .S1(net411),
    .X(_07194_));
 sky130_fd_sc_hd__mux4_2 _18839_ (.A0(_07190_),
    .A1(_07192_),
    .A2(_07193_),
    .A3(_07194_),
    .S0(net398),
    .S1(net396),
    .X(_07195_));
 sky130_fd_sc_hd__mux2i_4 _18840_ (.A0(_07189_),
    .A1(_07195_),
    .S(net394),
    .Y(_11593_));
 sky130_fd_sc_hd__mux4_2 _18841_ (.A0(\w[1][3] ),
    .A1(\w[5][3] ),
    .A2(\w[3][3] ),
    .A3(\w[7][3] ),
    .S0(net405),
    .S1(net409),
    .X(_07196_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1095 ();
 sky130_fd_sc_hd__mux4_2 _18843_ (.A0(\w[9][3] ),
    .A1(\w[13][3] ),
    .A2(\w[11][3] ),
    .A3(\w[15][3] ),
    .S0(net405),
    .S1(net409),
    .X(_07198_));
 sky130_fd_sc_hd__mux4_2 _18844_ (.A0(\w[17][3] ),
    .A1(\w[21][3] ),
    .A2(\w[19][3] ),
    .A3(\w[23][3] ),
    .S0(net405),
    .S1(net409),
    .X(_07199_));
 sky130_fd_sc_hd__mux4_2 _18845_ (.A0(\w[25][3] ),
    .A1(\w[29][3] ),
    .A2(\w[27][3] ),
    .A3(\w[31][3] ),
    .S0(net405),
    .S1(net409),
    .X(_07200_));
 sky130_fd_sc_hd__mux4_2 _18846_ (.A0(_07196_),
    .A1(_07198_),
    .A2(_07199_),
    .A3(_07200_),
    .S0(net400),
    .S1(net536),
    .X(_07201_));
 sky130_fd_sc_hd__mux4_2 _18847_ (.A0(\w[33][3] ),
    .A1(\w[37][3] ),
    .A2(\w[35][3] ),
    .A3(\w[39][3] ),
    .S0(net405),
    .S1(net409),
    .X(_07202_));
 sky130_fd_sc_hd__mux4_2 _18848_ (.A0(\w[41][3] ),
    .A1(\w[45][3] ),
    .A2(\w[43][3] ),
    .A3(\w[47][3] ),
    .S0(net405),
    .S1(net409),
    .X(_07203_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1094 ();
 sky130_fd_sc_hd__mux4_2 _18850_ (.A0(\w[49][3] ),
    .A1(\w[53][3] ),
    .A2(\w[51][3] ),
    .A3(\w[55][3] ),
    .S0(net405),
    .S1(net409),
    .X(_07205_));
 sky130_fd_sc_hd__mux4_2 _18851_ (.A0(\w[57][3] ),
    .A1(\w[61][3] ),
    .A2(\w[59][3] ),
    .A3(\w[63][3] ),
    .S0(net405),
    .S1(net409),
    .X(_07206_));
 sky130_fd_sc_hd__mux4_2 _18852_ (.A0(_07202_),
    .A1(_07203_),
    .A2(_07205_),
    .A3(_07206_),
    .S0(net400),
    .S1(net536),
    .X(_07207_));
 sky130_fd_sc_hd__mux2i_4 _18853_ (.A0(_07201_),
    .A1(_07207_),
    .S(net395),
    .Y(_11604_));
 sky130_fd_sc_hd__mux4_2 _18854_ (.A0(\w[1][4] ),
    .A1(\w[5][4] ),
    .A2(\w[3][4] ),
    .A3(\w[7][4] ),
    .S0(net401),
    .S1(net408),
    .X(_07208_));
 sky130_fd_sc_hd__mux4_2 _18855_ (.A0(\w[9][4] ),
    .A1(\w[13][4] ),
    .A2(\w[11][4] ),
    .A3(\w[15][4] ),
    .S0(net401),
    .S1(net408),
    .X(_07209_));
 sky130_fd_sc_hd__mux4_2 _18856_ (.A0(\w[17][4] ),
    .A1(\w[21][4] ),
    .A2(\w[19][4] ),
    .A3(\w[23][4] ),
    .S0(net401),
    .S1(net408),
    .X(_07210_));
 sky130_fd_sc_hd__mux4_2 _18857_ (.A0(\w[25][4] ),
    .A1(\w[29][4] ),
    .A2(\w[27][4] ),
    .A3(\w[31][4] ),
    .S0(net401),
    .S1(net408),
    .X(_07211_));
 sky130_fd_sc_hd__mux4_2 _18858_ (.A0(_07208_),
    .A1(_07209_),
    .A2(_07210_),
    .A3(_07211_),
    .S0(net398),
    .S1(net396),
    .X(_07212_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1093 ();
 sky130_fd_sc_hd__mux4_2 _18860_ (.A0(\w[33][4] ),
    .A1(\w[37][4] ),
    .A2(\w[35][4] ),
    .A3(\w[39][4] ),
    .S0(net404),
    .S1(net411),
    .X(_07214_));
 sky130_fd_sc_hd__mux4_2 _18861_ (.A0(\w[41][4] ),
    .A1(\w[45][4] ),
    .A2(\w[43][4] ),
    .A3(\w[47][4] ),
    .S0(net404),
    .S1(net411),
    .X(_07215_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1092 ();
 sky130_fd_sc_hd__mux4_2 _18863_ (.A0(\w[49][4] ),
    .A1(\w[53][4] ),
    .A2(\w[51][4] ),
    .A3(\w[55][4] ),
    .S0(net404),
    .S1(net411),
    .X(_07217_));
 sky130_fd_sc_hd__mux4_2 _18864_ (.A0(\w[57][4] ),
    .A1(\w[61][4] ),
    .A2(\w[59][4] ),
    .A3(\w[63][4] ),
    .S0(net404),
    .S1(net411),
    .X(_07218_));
 sky130_fd_sc_hd__mux4_2 _18865_ (.A0(_07214_),
    .A1(_07215_),
    .A2(_07217_),
    .A3(_07218_),
    .S0(net398),
    .S1(net396),
    .X(_07219_));
 sky130_fd_sc_hd__mux2i_4 _18866_ (.A0(_07212_),
    .A1(_07219_),
    .S(net394),
    .Y(_11612_));
 sky130_fd_sc_hd__mux4_2 _18867_ (.A0(\w[1][5] ),
    .A1(\w[5][5] ),
    .A2(\w[3][5] ),
    .A3(\w[7][5] ),
    .S0(net405),
    .S1(net409),
    .X(_07220_));
 sky130_fd_sc_hd__mux4_2 _18868_ (.A0(\w[9][5] ),
    .A1(\w[13][5] ),
    .A2(\w[11][5] ),
    .A3(\w[15][5] ),
    .S0(net405),
    .S1(net409),
    .X(_07221_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1091 ();
 sky130_fd_sc_hd__mux4_2 _18870_ (.A0(\w[17][5] ),
    .A1(\w[21][5] ),
    .A2(\w[19][5] ),
    .A3(\w[23][5] ),
    .S0(net405),
    .S1(net409),
    .X(_07223_));
 sky130_fd_sc_hd__mux4_2 _18871_ (.A0(\w[25][5] ),
    .A1(\w[29][5] ),
    .A2(\w[27][5] ),
    .A3(\w[31][5] ),
    .S0(net405),
    .S1(net409),
    .X(_07224_));
 sky130_fd_sc_hd__mux4_2 _18872_ (.A0(_07220_),
    .A1(_07221_),
    .A2(_07223_),
    .A3(_07224_),
    .S0(net400),
    .S1(net396),
    .X(_07225_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1090 ();
 sky130_fd_sc_hd__mux4_2 _18874_ (.A0(\w[33][5] ),
    .A1(\w[37][5] ),
    .A2(\w[35][5] ),
    .A3(\w[39][5] ),
    .S0(net405),
    .S1(net409),
    .X(_07227_));
 sky130_fd_sc_hd__mux4_2 _18875_ (.A0(\w[41][5] ),
    .A1(\w[45][5] ),
    .A2(\w[43][5] ),
    .A3(\w[47][5] ),
    .S0(net405),
    .S1(net409),
    .X(_07228_));
 sky130_fd_sc_hd__mux4_2 _18876_ (.A0(\w[49][5] ),
    .A1(\w[53][5] ),
    .A2(\w[51][5] ),
    .A3(\w[55][5] ),
    .S0(net405),
    .S1(net409),
    .X(_07229_));
 sky130_fd_sc_hd__mux4_2 _18877_ (.A0(\w[57][5] ),
    .A1(\w[61][5] ),
    .A2(\w[59][5] ),
    .A3(\w[63][5] ),
    .S0(net405),
    .S1(net409),
    .X(_07230_));
 sky130_fd_sc_hd__mux4_2 _18878_ (.A0(_07227_),
    .A1(_07228_),
    .A2(_07229_),
    .A3(_07230_),
    .S0(net400),
    .S1(net536),
    .X(_07231_));
 sky130_fd_sc_hd__mux2i_4 _18879_ (.A0(_07225_),
    .A1(_07231_),
    .S(net395),
    .Y(_11620_));
 sky130_fd_sc_hd__mux4_2 _18880_ (.A0(\w[1][6] ),
    .A1(\w[5][6] ),
    .A2(\w[3][6] ),
    .A3(\w[7][6] ),
    .S0(net403),
    .S1(net411),
    .X(_07232_));
 sky130_fd_sc_hd__mux4_2 _18881_ (.A0(\w[9][6] ),
    .A1(\w[13][6] ),
    .A2(\w[11][6] ),
    .A3(\w[15][6] ),
    .S0(net403),
    .S1(net411),
    .X(_07233_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1089 ();
 sky130_fd_sc_hd__mux4_2 _18883_ (.A0(\w[17][6] ),
    .A1(\w[21][6] ),
    .A2(\w[19][6] ),
    .A3(\w[23][6] ),
    .S0(net403),
    .S1(net411),
    .X(_07235_));
 sky130_fd_sc_hd__mux4_2 _18884_ (.A0(\w[25][6] ),
    .A1(\w[29][6] ),
    .A2(\w[27][6] ),
    .A3(\w[31][6] ),
    .S0(net403),
    .S1(net411),
    .X(_07236_));
 sky130_fd_sc_hd__mux4_2 _18885_ (.A0(_07232_),
    .A1(_07233_),
    .A2(_07235_),
    .A3(_07236_),
    .S0(net398),
    .S1(net396),
    .X(_07237_));
 sky130_fd_sc_hd__mux4_2 _18886_ (.A0(\w[33][6] ),
    .A1(\w[37][6] ),
    .A2(\w[35][6] ),
    .A3(\w[39][6] ),
    .S0(net404),
    .S1(net410),
    .X(_07238_));
 sky130_fd_sc_hd__mux4_2 _18887_ (.A0(\w[41][6] ),
    .A1(\w[45][6] ),
    .A2(\w[43][6] ),
    .A3(\w[47][6] ),
    .S0(net404),
    .S1(net410),
    .X(_07239_));
 sky130_fd_sc_hd__mux4_2 _18888_ (.A0(\w[49][6] ),
    .A1(\w[53][6] ),
    .A2(\w[51][6] ),
    .A3(\w[55][6] ),
    .S0(net404),
    .S1(net410),
    .X(_07240_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1088 ();
 sky130_fd_sc_hd__mux4_2 _18890_ (.A0(\w[57][6] ),
    .A1(\w[61][6] ),
    .A2(\w[59][6] ),
    .A3(\w[63][6] ),
    .S0(net404),
    .S1(net410),
    .X(_07242_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1087 ();
 sky130_fd_sc_hd__mux4_2 _18892_ (.A0(_07238_),
    .A1(_07239_),
    .A2(_07240_),
    .A3(_07242_),
    .S0(net537),
    .S1(net396),
    .X(_07244_));
 sky130_fd_sc_hd__mux2i_4 _18893_ (.A0(_07237_),
    .A1(_07244_),
    .S(net394),
    .Y(_11628_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1086 ();
 sky130_fd_sc_hd__mux4_2 _18895_ (.A0(\w[1][7] ),
    .A1(\w[5][7] ),
    .A2(\w[3][7] ),
    .A3(\w[7][7] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07246_));
 sky130_fd_sc_hd__mux4_2 _18896_ (.A0(\w[9][7] ),
    .A1(\w[13][7] ),
    .A2(\w[11][7] ),
    .A3(\w[15][7] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07247_));
 sky130_fd_sc_hd__mux4_2 _18897_ (.A0(\w[17][7] ),
    .A1(\w[21][7] ),
    .A2(\w[19][7] ),
    .A3(\w[23][7] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07248_));
 sky130_fd_sc_hd__mux4_2 _18898_ (.A0(\w[25][7] ),
    .A1(\w[29][7] ),
    .A2(\w[27][7] ),
    .A3(\w[31][7] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07249_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1085 ();
 sky130_fd_sc_hd__mux4_2 _18900_ (.A0(_07246_),
    .A1(_07247_),
    .A2(_07248_),
    .A3(_07249_),
    .S0(net400),
    .S1(\count7_1[4] ),
    .X(_07251_));
 sky130_fd_sc_hd__mux4_2 _18901_ (.A0(\w[33][7] ),
    .A1(\w[37][7] ),
    .A2(\w[35][7] ),
    .A3(\w[39][7] ),
    .S0(net405),
    .S1(net409),
    .X(_07252_));
 sky130_fd_sc_hd__mux4_2 _18902_ (.A0(\w[41][7] ),
    .A1(\w[45][7] ),
    .A2(\w[43][7] ),
    .A3(\w[47][7] ),
    .S0(net405),
    .S1(net409),
    .X(_07253_));
 sky130_fd_sc_hd__mux4_2 _18903_ (.A0(\w[49][7] ),
    .A1(\w[53][7] ),
    .A2(\w[51][7] ),
    .A3(\w[55][7] ),
    .S0(net405),
    .S1(net409),
    .X(_07254_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1084 ();
 sky130_fd_sc_hd__mux4_2 _18905_ (.A0(\w[57][7] ),
    .A1(\w[61][7] ),
    .A2(\w[59][7] ),
    .A3(\w[63][7] ),
    .S0(net405),
    .S1(net409),
    .X(_07256_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1083 ();
 sky130_fd_sc_hd__mux4_2 _18907_ (.A0(_07252_),
    .A1(_07253_),
    .A2(_07254_),
    .A3(_07256_),
    .S0(net400),
    .S1(net536),
    .X(_07258_));
 sky130_fd_sc_hd__mux2i_4 _18908_ (.A0(_07251_),
    .A1(_07258_),
    .S(net395),
    .Y(_11636_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1082 ();
 sky130_fd_sc_hd__mux4_2 _18910_ (.A0(\w[1][8] ),
    .A1(\w[5][8] ),
    .A2(\w[3][8] ),
    .A3(\w[7][8] ),
    .S0(net403),
    .S1(net411),
    .X(_07260_));
 sky130_fd_sc_hd__mux4_2 _18911_ (.A0(\w[9][8] ),
    .A1(\w[13][8] ),
    .A2(\w[11][8] ),
    .A3(\w[15][8] ),
    .S0(net403),
    .S1(net411),
    .X(_07261_));
 sky130_fd_sc_hd__mux4_2 _18912_ (.A0(\w[17][8] ),
    .A1(\w[21][8] ),
    .A2(\w[19][8] ),
    .A3(\w[23][8] ),
    .S0(net403),
    .S1(net411),
    .X(_07262_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1081 ();
 sky130_fd_sc_hd__mux4_2 _18914_ (.A0(\w[25][8] ),
    .A1(\w[29][8] ),
    .A2(\w[27][8] ),
    .A3(\w[31][8] ),
    .S0(net403),
    .S1(net411),
    .X(_07264_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1080 ();
 sky130_fd_sc_hd__mux4_2 _18916_ (.A0(_07260_),
    .A1(_07261_),
    .A2(_07262_),
    .A3(_07264_),
    .S0(net398),
    .S1(net396),
    .X(_07266_));
 sky130_fd_sc_hd__mux4_2 _18917_ (.A0(\w[33][8] ),
    .A1(\w[37][8] ),
    .A2(\w[35][8] ),
    .A3(\w[39][8] ),
    .S0(net404),
    .S1(net410),
    .X(_07267_));
 sky130_fd_sc_hd__mux4_2 _18918_ (.A0(\w[41][8] ),
    .A1(\w[45][8] ),
    .A2(\w[43][8] ),
    .A3(\w[47][8] ),
    .S0(net404),
    .S1(net410),
    .X(_07268_));
 sky130_fd_sc_hd__mux4_2 _18919_ (.A0(\w[49][8] ),
    .A1(\w[53][8] ),
    .A2(\w[51][8] ),
    .A3(\w[55][8] ),
    .S0(net404),
    .S1(net410),
    .X(_07269_));
 sky130_fd_sc_hd__mux4_2 _18920_ (.A0(\w[57][8] ),
    .A1(\w[61][8] ),
    .A2(\w[59][8] ),
    .A3(\w[63][8] ),
    .S0(net404),
    .S1(net410),
    .X(_07270_));
 sky130_fd_sc_hd__mux4_2 _18921_ (.A0(_07267_),
    .A1(_07268_),
    .A2(_07269_),
    .A3(_07270_),
    .S0(net537),
    .S1(net397),
    .X(_07271_));
 sky130_fd_sc_hd__mux2i_4 _18922_ (.A0(_07266_),
    .A1(_07271_),
    .S(net394),
    .Y(_11644_));
 sky130_fd_sc_hd__mux4_2 _18923_ (.A0(\w[1][9] ),
    .A1(\w[5][9] ),
    .A2(\w[3][9] ),
    .A3(\w[7][9] ),
    .S0(net407),
    .S1(net409),
    .X(_07272_));
 sky130_fd_sc_hd__mux4_2 _18924_ (.A0(\w[9][9] ),
    .A1(\w[13][9] ),
    .A2(\w[11][9] ),
    .A3(\w[15][9] ),
    .S0(net407),
    .S1(net409),
    .X(_07273_));
 sky130_fd_sc_hd__mux4_2 _18925_ (.A0(\w[17][9] ),
    .A1(\w[21][9] ),
    .A2(\w[19][9] ),
    .A3(\w[23][9] ),
    .S0(net407),
    .S1(net409),
    .X(_07274_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1079 ();
 sky130_fd_sc_hd__mux4_2 _18927_ (.A0(\w[25][9] ),
    .A1(\w[29][9] ),
    .A2(\w[27][9] ),
    .A3(\w[31][9] ),
    .S0(net407),
    .S1(net409),
    .X(_07276_));
 sky130_fd_sc_hd__mux4_2 _18928_ (.A0(_07272_),
    .A1(_07273_),
    .A2(_07274_),
    .A3(_07276_),
    .S0(net400),
    .S1(\count7_1[4] ),
    .X(_07277_));
 sky130_fd_sc_hd__mux4_2 _18929_ (.A0(\w[33][9] ),
    .A1(\w[37][9] ),
    .A2(\w[35][9] ),
    .A3(\w[39][9] ),
    .S0(net406),
    .S1(net412),
    .X(_07278_));
 sky130_fd_sc_hd__mux4_2 _18930_ (.A0(\w[41][9] ),
    .A1(\w[45][9] ),
    .A2(\w[43][9] ),
    .A3(\w[47][9] ),
    .S0(net406),
    .S1(net412),
    .X(_07279_));
 sky130_fd_sc_hd__mux4_2 _18931_ (.A0(\w[49][9] ),
    .A1(\w[53][9] ),
    .A2(\w[51][9] ),
    .A3(\w[55][9] ),
    .S0(net406),
    .S1(net412),
    .X(_07280_));
 sky130_fd_sc_hd__mux4_2 _18932_ (.A0(\w[57][9] ),
    .A1(\w[61][9] ),
    .A2(\w[59][9] ),
    .A3(\w[63][9] ),
    .S0(net406),
    .S1(net412),
    .X(_07281_));
 sky130_fd_sc_hd__mux4_2 _18933_ (.A0(_07278_),
    .A1(_07279_),
    .A2(_07280_),
    .A3(_07281_),
    .S0(net537),
    .S1(net396),
    .X(_07282_));
 sky130_fd_sc_hd__mux2i_4 _18934_ (.A0(_07277_),
    .A1(_07282_),
    .S(\count7_1[5] ),
    .Y(_11652_));
 sky130_fd_sc_hd__mux4_2 _18935_ (.A0(\w[1][10] ),
    .A1(\w[5][10] ),
    .A2(\w[3][10] ),
    .A3(\w[7][10] ),
    .S0(net402),
    .S1(net410),
    .X(_07283_));
 sky130_fd_sc_hd__mux4_2 _18936_ (.A0(\w[9][10] ),
    .A1(\w[13][10] ),
    .A2(\w[11][10] ),
    .A3(\w[15][10] ),
    .S0(net402),
    .S1(net410),
    .X(_07284_));
 sky130_fd_sc_hd__mux4_2 _18937_ (.A0(\w[17][10] ),
    .A1(\w[21][10] ),
    .A2(\w[19][10] ),
    .A3(\w[23][10] ),
    .S0(net402),
    .S1(net410),
    .X(_07285_));
 sky130_fd_sc_hd__mux4_2 _18938_ (.A0(\w[25][10] ),
    .A1(\w[29][10] ),
    .A2(\w[27][10] ),
    .A3(\w[31][10] ),
    .S0(net402),
    .S1(net410),
    .X(_07286_));
 sky130_fd_sc_hd__mux4_2 _18939_ (.A0(_07283_),
    .A1(_07284_),
    .A2(_07285_),
    .A3(_07286_),
    .S0(net399),
    .S1(net397),
    .X(_07287_));
 sky130_fd_sc_hd__mux4_2 _18940_ (.A0(\w[33][10] ),
    .A1(\w[37][10] ),
    .A2(\w[35][10] ),
    .A3(\w[39][10] ),
    .S0(net402),
    .S1(net410),
    .X(_07288_));
 sky130_fd_sc_hd__mux4_2 _18941_ (.A0(\w[41][10] ),
    .A1(\w[45][10] ),
    .A2(\w[43][10] ),
    .A3(\w[47][10] ),
    .S0(net402),
    .S1(net410),
    .X(_07289_));
 sky130_fd_sc_hd__mux4_2 _18942_ (.A0(\w[49][10] ),
    .A1(\w[53][10] ),
    .A2(\w[51][10] ),
    .A3(\w[55][10] ),
    .S0(net402),
    .S1(net410),
    .X(_07290_));
 sky130_fd_sc_hd__mux4_2 _18943_ (.A0(\w[57][10] ),
    .A1(\w[61][10] ),
    .A2(\w[59][10] ),
    .A3(\w[63][10] ),
    .S0(net402),
    .S1(net410),
    .X(_07291_));
 sky130_fd_sc_hd__mux4_2 _18944_ (.A0(_07288_),
    .A1(_07289_),
    .A2(_07290_),
    .A3(_07291_),
    .S0(net399),
    .S1(net397),
    .X(_07292_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1078 ();
 sky130_fd_sc_hd__mux2i_4 _18946_ (.A0(_07287_),
    .A1(_07292_),
    .S(net394),
    .Y(_11660_));
 sky130_fd_sc_hd__mux4_2 _18947_ (.A0(\w[1][11] ),
    .A1(\w[5][11] ),
    .A2(\w[3][11] ),
    .A3(\w[7][11] ),
    .S0(net403),
    .S1(net411),
    .X(_07294_));
 sky130_fd_sc_hd__mux4_2 _18948_ (.A0(\w[9][11] ),
    .A1(\w[13][11] ),
    .A2(\w[11][11] ),
    .A3(\w[15][11] ),
    .S0(net403),
    .S1(net411),
    .X(_07295_));
 sky130_fd_sc_hd__mux4_2 _18949_ (.A0(\w[17][11] ),
    .A1(\w[21][11] ),
    .A2(\w[19][11] ),
    .A3(\w[23][11] ),
    .S0(net403),
    .S1(net411),
    .X(_07296_));
 sky130_fd_sc_hd__mux4_2 _18950_ (.A0(\w[25][11] ),
    .A1(\w[29][11] ),
    .A2(\w[27][11] ),
    .A3(\w[31][11] ),
    .S0(net403),
    .S1(net411),
    .X(_07297_));
 sky130_fd_sc_hd__mux4_2 _18951_ (.A0(_07294_),
    .A1(_07295_),
    .A2(_07296_),
    .A3(_07297_),
    .S0(net398),
    .S1(net396),
    .X(_07298_));
 sky130_fd_sc_hd__mux4_2 _18952_ (.A0(\w[33][11] ),
    .A1(\w[37][11] ),
    .A2(\w[35][11] ),
    .A3(\w[39][11] ),
    .S0(net538),
    .S1(net412),
    .X(_07299_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1077 ();
 sky130_fd_sc_hd__mux4_2 _18954_ (.A0(\w[41][11] ),
    .A1(\w[45][11] ),
    .A2(\w[43][11] ),
    .A3(\w[47][11] ),
    .S0(net538),
    .S1(net412),
    .X(_07301_));
 sky130_fd_sc_hd__mux4_2 _18955_ (.A0(\w[49][11] ),
    .A1(\w[53][11] ),
    .A2(\w[51][11] ),
    .A3(\w[55][11] ),
    .S0(net538),
    .S1(net412),
    .X(_07302_));
 sky130_fd_sc_hd__mux4_2 _18956_ (.A0(\w[57][11] ),
    .A1(\w[61][11] ),
    .A2(\w[59][11] ),
    .A3(\w[63][11] ),
    .S0(net538),
    .S1(net412),
    .X(_07303_));
 sky130_fd_sc_hd__mux4_2 _18957_ (.A0(_07299_),
    .A1(_07301_),
    .A2(_07302_),
    .A3(_07303_),
    .S0(net399),
    .S1(net397),
    .X(_07304_));
 sky130_fd_sc_hd__mux2i_2 _18958_ (.A0(_07298_),
    .A1(_07304_),
    .S(\count7_1[5] ),
    .Y(_11668_));
 sky130_fd_sc_hd__mux4_2 _18959_ (.A0(\w[1][12] ),
    .A1(\w[5][12] ),
    .A2(\w[3][12] ),
    .A3(\w[7][12] ),
    .S0(net403),
    .S1(net411),
    .X(_07305_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1076 ();
 sky130_fd_sc_hd__mux4_2 _18961_ (.A0(\w[9][12] ),
    .A1(\w[13][12] ),
    .A2(\w[11][12] ),
    .A3(\w[15][12] ),
    .S0(net403),
    .S1(net411),
    .X(_07307_));
 sky130_fd_sc_hd__mux4_2 _18962_ (.A0(\w[17][12] ),
    .A1(\w[21][12] ),
    .A2(\w[19][12] ),
    .A3(\w[23][12] ),
    .S0(net403),
    .S1(net411),
    .X(_07308_));
 sky130_fd_sc_hd__mux4_2 _18963_ (.A0(\w[25][12] ),
    .A1(\w[29][12] ),
    .A2(\w[27][12] ),
    .A3(\w[31][12] ),
    .S0(net403),
    .S1(net411),
    .X(_07309_));
 sky130_fd_sc_hd__mux4_2 _18964_ (.A0(_07305_),
    .A1(_07307_),
    .A2(_07308_),
    .A3(_07309_),
    .S0(net399),
    .S1(net397),
    .X(_07310_));
 sky130_fd_sc_hd__mux4_2 _18965_ (.A0(\w[33][12] ),
    .A1(\w[37][12] ),
    .A2(\w[35][12] ),
    .A3(\w[39][12] ),
    .S0(net402),
    .S1(net410),
    .X(_07311_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1075 ();
 sky130_fd_sc_hd__mux4_2 _18967_ (.A0(\w[41][12] ),
    .A1(\w[45][12] ),
    .A2(\w[43][12] ),
    .A3(\w[47][12] ),
    .S0(net402),
    .S1(net410),
    .X(_07313_));
 sky130_fd_sc_hd__mux4_2 _18968_ (.A0(\w[49][12] ),
    .A1(\w[53][12] ),
    .A2(\w[51][12] ),
    .A3(\w[55][12] ),
    .S0(net402),
    .S1(net410),
    .X(_07314_));
 sky130_fd_sc_hd__mux4_2 _18969_ (.A0(\w[57][12] ),
    .A1(\w[61][12] ),
    .A2(\w[59][12] ),
    .A3(\w[63][12] ),
    .S0(net402),
    .S1(net410),
    .X(_07315_));
 sky130_fd_sc_hd__mux4_2 _18970_ (.A0(_07311_),
    .A1(_07313_),
    .A2(_07314_),
    .A3(_07315_),
    .S0(net399),
    .S1(net397),
    .X(_07316_));
 sky130_fd_sc_hd__mux2i_4 _18971_ (.A0(_07310_),
    .A1(_07316_),
    .S(net394),
    .Y(_11676_));
 sky130_fd_sc_hd__mux4_2 _18972_ (.A0(\w[1][13] ),
    .A1(\w[5][13] ),
    .A2(\w[3][13] ),
    .A3(\w[7][13] ),
    .S0(net402),
    .S1(net410),
    .X(_07317_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1074 ();
 sky130_fd_sc_hd__mux4_2 _18974_ (.A0(\w[9][13] ),
    .A1(\w[13][13] ),
    .A2(\w[11][13] ),
    .A3(\w[15][13] ),
    .S0(net402),
    .S1(net410),
    .X(_07319_));
 sky130_fd_sc_hd__mux4_2 _18975_ (.A0(\w[17][13] ),
    .A1(\w[21][13] ),
    .A2(\w[19][13] ),
    .A3(\w[23][13] ),
    .S0(net402),
    .S1(net410),
    .X(_07320_));
 sky130_fd_sc_hd__mux4_2 _18976_ (.A0(\w[25][13] ),
    .A1(\w[29][13] ),
    .A2(\w[27][13] ),
    .A3(\w[31][13] ),
    .S0(net402),
    .S1(net410),
    .X(_07321_));
 sky130_fd_sc_hd__mux4_2 _18977_ (.A0(_07317_),
    .A1(_07319_),
    .A2(_07320_),
    .A3(_07321_),
    .S0(net399),
    .S1(net397),
    .X(_07322_));
 sky130_fd_sc_hd__mux4_2 _18978_ (.A0(\w[33][13] ),
    .A1(\w[37][13] ),
    .A2(\w[35][13] ),
    .A3(\w[39][13] ),
    .S0(net538),
    .S1(net412),
    .X(_07323_));
 sky130_fd_sc_hd__mux4_2 _18979_ (.A0(\w[41][13] ),
    .A1(\w[45][13] ),
    .A2(\w[43][13] ),
    .A3(\w[47][13] ),
    .S0(net538),
    .S1(net412),
    .X(_07324_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1073 ();
 sky130_fd_sc_hd__mux4_2 _18981_ (.A0(\w[49][13] ),
    .A1(\w[53][13] ),
    .A2(\w[51][13] ),
    .A3(\w[55][13] ),
    .S0(net538),
    .S1(net412),
    .X(_07326_));
 sky130_fd_sc_hd__mux4_2 _18982_ (.A0(\w[57][13] ),
    .A1(\w[61][13] ),
    .A2(\w[59][13] ),
    .A3(\w[63][13] ),
    .S0(net538),
    .S1(net412),
    .X(_07327_));
 sky130_fd_sc_hd__mux4_2 _18983_ (.A0(_07323_),
    .A1(_07324_),
    .A2(_07326_),
    .A3(_07327_),
    .S0(net399),
    .S1(net397),
    .X(_07328_));
 sky130_fd_sc_hd__mux2i_4 _18984_ (.A0(_07322_),
    .A1(_07328_),
    .S(\count7_1[5] ),
    .Y(_11684_));
 sky130_fd_sc_hd__mux4_2 _18985_ (.A0(\w[1][14] ),
    .A1(\w[5][14] ),
    .A2(\w[3][14] ),
    .A3(\w[7][14] ),
    .S0(net404),
    .S1(net408),
    .X(_07329_));
 sky130_fd_sc_hd__mux4_2 _18986_ (.A0(\w[9][14] ),
    .A1(\w[13][14] ),
    .A2(\w[11][14] ),
    .A3(\w[15][14] ),
    .S0(net404),
    .S1(net408),
    .X(_07330_));
 sky130_fd_sc_hd__mux4_2 _18987_ (.A0(\w[17][14] ),
    .A1(\w[21][14] ),
    .A2(\w[19][14] ),
    .A3(\w[23][14] ),
    .S0(net404),
    .S1(net408),
    .X(_07331_));
 sky130_fd_sc_hd__mux4_2 _18988_ (.A0(\w[25][14] ),
    .A1(\w[29][14] ),
    .A2(\w[27][14] ),
    .A3(\w[31][14] ),
    .S0(net404),
    .S1(net408),
    .X(_07332_));
 sky130_fd_sc_hd__mux4_2 _18989_ (.A0(_07329_),
    .A1(_07330_),
    .A2(_07331_),
    .A3(_07332_),
    .S0(net398),
    .S1(net396),
    .X(_07333_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1072 ();
 sky130_fd_sc_hd__mux4_2 _18991_ (.A0(\w[33][14] ),
    .A1(\w[37][14] ),
    .A2(\w[35][14] ),
    .A3(\w[39][14] ),
    .S0(net403),
    .S1(net411),
    .X(_07335_));
 sky130_fd_sc_hd__mux4_2 _18992_ (.A0(\w[41][14] ),
    .A1(\w[45][14] ),
    .A2(\w[43][14] ),
    .A3(\w[47][14] ),
    .S0(net403),
    .S1(net411),
    .X(_07336_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1071 ();
 sky130_fd_sc_hd__mux4_2 _18994_ (.A0(\w[49][14] ),
    .A1(\w[53][14] ),
    .A2(\w[51][14] ),
    .A3(\w[55][14] ),
    .S0(net403),
    .S1(net411),
    .X(_07338_));
 sky130_fd_sc_hd__mux4_2 _18995_ (.A0(\w[57][14] ),
    .A1(\w[61][14] ),
    .A2(\w[59][14] ),
    .A3(\w[63][14] ),
    .S0(net403),
    .S1(net411),
    .X(_07339_));
 sky130_fd_sc_hd__mux4_2 _18996_ (.A0(_07335_),
    .A1(_07336_),
    .A2(_07338_),
    .A3(_07339_),
    .S0(net537),
    .S1(net396),
    .X(_07340_));
 sky130_fd_sc_hd__mux2i_4 _18997_ (.A0(_07333_),
    .A1(_07340_),
    .S(net394),
    .Y(_11692_));
 sky130_fd_sc_hd__mux4_2 _18998_ (.A0(\w[1][15] ),
    .A1(\w[5][15] ),
    .A2(\w[3][15] ),
    .A3(\w[7][15] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07341_));
 sky130_fd_sc_hd__mux4_2 _18999_ (.A0(\w[9][15] ),
    .A1(\w[13][15] ),
    .A2(\w[11][15] ),
    .A3(\w[15][15] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07342_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1070 ();
 sky130_fd_sc_hd__mux4_2 _19001_ (.A0(\w[17][15] ),
    .A1(\w[21][15] ),
    .A2(\w[19][15] ),
    .A3(\w[23][15] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07344_));
 sky130_fd_sc_hd__mux4_2 _19002_ (.A0(\w[25][15] ),
    .A1(\w[29][15] ),
    .A2(\w[27][15] ),
    .A3(\w[31][15] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07345_));
 sky130_fd_sc_hd__mux4_2 _19003_ (.A0(_07341_),
    .A1(_07342_),
    .A2(_07344_),
    .A3(_07345_),
    .S0(net400),
    .S1(\count7_1[4] ),
    .X(_07346_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1069 ();
 sky130_fd_sc_hd__mux4_2 _19005_ (.A0(\w[33][15] ),
    .A1(\w[37][15] ),
    .A2(\w[35][15] ),
    .A3(\w[39][15] ),
    .S0(net406),
    .S1(net412),
    .X(_07348_));
 sky130_fd_sc_hd__mux4_2 _19006_ (.A0(\w[41][15] ),
    .A1(\w[45][15] ),
    .A2(\w[43][15] ),
    .A3(\w[47][15] ),
    .S0(net406),
    .S1(net412),
    .X(_07349_));
 sky130_fd_sc_hd__mux4_2 _19007_ (.A0(\w[49][15] ),
    .A1(\w[53][15] ),
    .A2(\w[51][15] ),
    .A3(\w[55][15] ),
    .S0(\count7_1[2] ),
    .S1(net412),
    .X(_07350_));
 sky130_fd_sc_hd__mux4_2 _19008_ (.A0(\w[57][15] ),
    .A1(\w[61][15] ),
    .A2(\w[59][15] ),
    .A3(\w[63][15] ),
    .S0(\count7_1[2] ),
    .S1(net412),
    .X(_07351_));
 sky130_fd_sc_hd__mux4_2 _19009_ (.A0(_07348_),
    .A1(_07349_),
    .A2(_07350_),
    .A3(_07351_),
    .S0(net537),
    .S1(\count7_1[4] ),
    .X(_07352_));
 sky130_fd_sc_hd__mux2i_2 _19010_ (.A0(_07346_),
    .A1(_07352_),
    .S(\count7_1[5] ),
    .Y(_11700_));
 sky130_fd_sc_hd__mux4_2 _19011_ (.A0(\w[1][16] ),
    .A1(\w[5][16] ),
    .A2(\w[3][16] ),
    .A3(\w[7][16] ),
    .S0(net404),
    .S1(net408),
    .X(_07353_));
 sky130_fd_sc_hd__mux4_2 _19012_ (.A0(\w[9][16] ),
    .A1(\w[13][16] ),
    .A2(\w[11][16] ),
    .A3(\w[15][16] ),
    .S0(net404),
    .S1(net408),
    .X(_07354_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1068 ();
 sky130_fd_sc_hd__mux4_2 _19014_ (.A0(\w[17][16] ),
    .A1(\w[21][16] ),
    .A2(\w[19][16] ),
    .A3(\w[23][16] ),
    .S0(net404),
    .S1(net408),
    .X(_07356_));
 sky130_fd_sc_hd__mux4_2 _19015_ (.A0(\w[25][16] ),
    .A1(\w[29][16] ),
    .A2(\w[27][16] ),
    .A3(\w[31][16] ),
    .S0(net404),
    .S1(net408),
    .X(_07357_));
 sky130_fd_sc_hd__mux4_2 _19016_ (.A0(_07353_),
    .A1(_07354_),
    .A2(_07356_),
    .A3(_07357_),
    .S0(net398),
    .S1(net396),
    .X(_07358_));
 sky130_fd_sc_hd__mux4_2 _19017_ (.A0(\w[33][16] ),
    .A1(\w[37][16] ),
    .A2(\w[35][16] ),
    .A3(\w[39][16] ),
    .S0(net402),
    .S1(net410),
    .X(_07359_));
 sky130_fd_sc_hd__mux4_2 _19018_ (.A0(\w[41][16] ),
    .A1(\w[45][16] ),
    .A2(\w[43][16] ),
    .A3(\w[47][16] ),
    .S0(net404),
    .S1(net410),
    .X(_07360_));
 sky130_fd_sc_hd__mux4_2 _19019_ (.A0(\w[49][16] ),
    .A1(\w[53][16] ),
    .A2(\w[51][16] ),
    .A3(\w[55][16] ),
    .S0(net404),
    .S1(net410),
    .X(_07361_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1067 ();
 sky130_fd_sc_hd__mux4_2 _19021_ (.A0(\w[57][16] ),
    .A1(\w[61][16] ),
    .A2(\w[59][16] ),
    .A3(\w[63][16] ),
    .S0(net404),
    .S1(net410),
    .X(_07363_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1066 ();
 sky130_fd_sc_hd__mux4_2 _19023_ (.A0(_07359_),
    .A1(_07360_),
    .A2(_07361_),
    .A3(_07363_),
    .S0(net537),
    .S1(net396),
    .X(_07365_));
 sky130_fd_sc_hd__mux2i_4 _19024_ (.A0(_07358_),
    .A1(_07365_),
    .S(net394),
    .Y(_11708_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1065 ();
 sky130_fd_sc_hd__mux4_2 _19026_ (.A0(\w[1][17] ),
    .A1(\w[5][17] ),
    .A2(\w[3][17] ),
    .A3(\w[7][17] ),
    .S0(net401),
    .S1(net408),
    .X(_07367_));
 sky130_fd_sc_hd__mux4_2 _19027_ (.A0(\w[9][17] ),
    .A1(\w[13][17] ),
    .A2(\w[11][17] ),
    .A3(\w[15][17] ),
    .S0(net401),
    .S1(net408),
    .X(_07368_));
 sky130_fd_sc_hd__mux4_2 _19028_ (.A0(\w[17][17] ),
    .A1(\w[21][17] ),
    .A2(\w[19][17] ),
    .A3(\w[23][17] ),
    .S0(net401),
    .S1(net408),
    .X(_07369_));
 sky130_fd_sc_hd__mux4_2 _19029_ (.A0(\w[25][17] ),
    .A1(\w[29][17] ),
    .A2(\w[27][17] ),
    .A3(\w[31][17] ),
    .S0(net401),
    .S1(net408),
    .X(_07370_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1064 ();
 sky130_fd_sc_hd__mux4_2 _19031_ (.A0(_07367_),
    .A1(_07368_),
    .A2(_07369_),
    .A3(_07370_),
    .S0(net398),
    .S1(net396),
    .X(_07372_));
 sky130_fd_sc_hd__mux4_2 _19032_ (.A0(\w[33][17] ),
    .A1(\w[37][17] ),
    .A2(\w[35][17] ),
    .A3(\w[39][17] ),
    .S0(net401),
    .S1(net408),
    .X(_07373_));
 sky130_fd_sc_hd__mux4_2 _19033_ (.A0(\w[41][17] ),
    .A1(\w[45][17] ),
    .A2(\w[43][17] ),
    .A3(\w[47][17] ),
    .S0(net401),
    .S1(net408),
    .X(_07374_));
 sky130_fd_sc_hd__mux4_2 _19034_ (.A0(\w[49][17] ),
    .A1(\w[53][17] ),
    .A2(\w[51][17] ),
    .A3(\w[55][17] ),
    .S0(net401),
    .S1(net408),
    .X(_07375_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1063 ();
 sky130_fd_sc_hd__mux4_2 _19036_ (.A0(\w[57][17] ),
    .A1(\w[61][17] ),
    .A2(\w[59][17] ),
    .A3(\w[63][17] ),
    .S0(net401),
    .S1(net408),
    .X(_07377_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1062 ();
 sky130_fd_sc_hd__mux4_2 _19038_ (.A0(_07373_),
    .A1(_07374_),
    .A2(_07375_),
    .A3(_07377_),
    .S0(net398),
    .S1(net396),
    .X(_07379_));
 sky130_fd_sc_hd__mux2i_4 _19039_ (.A0(_07372_),
    .A1(_07379_),
    .S(net394),
    .Y(_11716_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1061 ();
 sky130_fd_sc_hd__mux4_2 _19041_ (.A0(\w[1][18] ),
    .A1(\w[5][18] ),
    .A2(\w[3][18] ),
    .A3(\w[7][18] ),
    .S0(net402),
    .S1(net410),
    .X(_07381_));
 sky130_fd_sc_hd__mux4_2 _19042_ (.A0(\w[9][18] ),
    .A1(\w[13][18] ),
    .A2(\w[11][18] ),
    .A3(\w[15][18] ),
    .S0(net402),
    .S1(net410),
    .X(_07382_));
 sky130_fd_sc_hd__mux4_2 _19043_ (.A0(\w[17][18] ),
    .A1(\w[21][18] ),
    .A2(\w[19][18] ),
    .A3(\w[23][18] ),
    .S0(net402),
    .S1(net410),
    .X(_07383_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1060 ();
 sky130_fd_sc_hd__mux4_2 _19045_ (.A0(\w[25][18] ),
    .A1(\w[29][18] ),
    .A2(\w[27][18] ),
    .A3(\w[31][18] ),
    .S0(net402),
    .S1(net410),
    .X(_07385_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1059 ();
 sky130_fd_sc_hd__mux4_2 _19047_ (.A0(_07381_),
    .A1(_07382_),
    .A2(_07383_),
    .A3(_07385_),
    .S0(net399),
    .S1(net397),
    .X(_07387_));
 sky130_fd_sc_hd__mux4_2 _19048_ (.A0(\w[33][18] ),
    .A1(\w[37][18] ),
    .A2(\w[35][18] ),
    .A3(\w[39][18] ),
    .S0(net402),
    .S1(net410),
    .X(_07388_));
 sky130_fd_sc_hd__mux4_2 _19049_ (.A0(\w[41][18] ),
    .A1(\w[45][18] ),
    .A2(\w[43][18] ),
    .A3(\w[47][18] ),
    .S0(net402),
    .S1(net410),
    .X(_07389_));
 sky130_fd_sc_hd__mux4_2 _19050_ (.A0(\w[49][18] ),
    .A1(\w[53][18] ),
    .A2(\w[51][18] ),
    .A3(\w[55][18] ),
    .S0(net402),
    .S1(net410),
    .X(_07390_));
 sky130_fd_sc_hd__mux4_2 _19051_ (.A0(\w[57][18] ),
    .A1(\w[61][18] ),
    .A2(\w[59][18] ),
    .A3(\w[63][18] ),
    .S0(net402),
    .S1(net410),
    .X(_07391_));
 sky130_fd_sc_hd__mux4_2 _19052_ (.A0(_07388_),
    .A1(_07389_),
    .A2(_07390_),
    .A3(_07391_),
    .S0(net399),
    .S1(net397),
    .X(_07392_));
 sky130_fd_sc_hd__mux2i_4 _19053_ (.A0(_07387_),
    .A1(_07392_),
    .S(net394),
    .Y(_11724_));
 sky130_fd_sc_hd__mux4_2 _19054_ (.A0(\w[1][19] ),
    .A1(\w[5][19] ),
    .A2(\w[3][19] ),
    .A3(\w[7][19] ),
    .S0(net402),
    .S1(net410),
    .X(_07393_));
 sky130_fd_sc_hd__mux4_2 _19055_ (.A0(\w[9][19] ),
    .A1(\w[13][19] ),
    .A2(\w[11][19] ),
    .A3(\w[15][19] ),
    .S0(net402),
    .S1(net410),
    .X(_07394_));
 sky130_fd_sc_hd__mux4_2 _19056_ (.A0(\w[17][19] ),
    .A1(\w[21][19] ),
    .A2(\w[19][19] ),
    .A3(\w[23][19] ),
    .S0(net402),
    .S1(net410),
    .X(_07395_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1058 ();
 sky130_fd_sc_hd__mux4_2 _19058_ (.A0(\w[25][19] ),
    .A1(\w[29][19] ),
    .A2(\w[27][19] ),
    .A3(\w[31][19] ),
    .S0(net402),
    .S1(net410),
    .X(_07397_));
 sky130_fd_sc_hd__mux4_2 _19059_ (.A0(_07393_),
    .A1(_07394_),
    .A2(_07395_),
    .A3(_07397_),
    .S0(net399),
    .S1(net397),
    .X(_07398_));
 sky130_fd_sc_hd__mux4_2 _19060_ (.A0(\w[33][19] ),
    .A1(\w[37][19] ),
    .A2(\w[35][19] ),
    .A3(\w[39][19] ),
    .S0(net538),
    .S1(net412),
    .X(_07399_));
 sky130_fd_sc_hd__mux4_2 _19061_ (.A0(\w[41][19] ),
    .A1(\w[45][19] ),
    .A2(\w[43][19] ),
    .A3(\w[47][19] ),
    .S0(net538),
    .S1(net412),
    .X(_07400_));
 sky130_fd_sc_hd__mux4_2 _19062_ (.A0(\w[49][19] ),
    .A1(\w[53][19] ),
    .A2(\w[51][19] ),
    .A3(\w[55][19] ),
    .S0(net538),
    .S1(net412),
    .X(_07401_));
 sky130_fd_sc_hd__mux4_2 _19063_ (.A0(\w[57][19] ),
    .A1(\w[61][19] ),
    .A2(\w[59][19] ),
    .A3(\w[63][19] ),
    .S0(net538),
    .S1(net412),
    .X(_07402_));
 sky130_fd_sc_hd__mux4_2 _19064_ (.A0(_07399_),
    .A1(_07400_),
    .A2(_07401_),
    .A3(_07402_),
    .S0(net399),
    .S1(net397),
    .X(_07403_));
 sky130_fd_sc_hd__mux2i_4 _19065_ (.A0(_07398_),
    .A1(_07403_),
    .S(\count7_1[5] ),
    .Y(_11732_));
 sky130_fd_sc_hd__mux4_2 _19066_ (.A0(\w[1][20] ),
    .A1(\w[5][20] ),
    .A2(\w[3][20] ),
    .A3(\w[7][20] ),
    .S0(net402),
    .S1(net410),
    .X(_07404_));
 sky130_fd_sc_hd__mux4_2 _19067_ (.A0(\w[9][20] ),
    .A1(\w[13][20] ),
    .A2(\w[11][20] ),
    .A3(\w[15][20] ),
    .S0(net402),
    .S1(net410),
    .X(_07405_));
 sky130_fd_sc_hd__mux4_2 _19068_ (.A0(\w[17][20] ),
    .A1(\w[21][20] ),
    .A2(\w[19][20] ),
    .A3(\w[23][20] ),
    .S0(net402),
    .S1(net410),
    .X(_07406_));
 sky130_fd_sc_hd__mux4_2 _19069_ (.A0(\w[25][20] ),
    .A1(\w[29][20] ),
    .A2(\w[27][20] ),
    .A3(\w[31][20] ),
    .S0(net402),
    .S1(net410),
    .X(_07407_));
 sky130_fd_sc_hd__mux4_2 _19070_ (.A0(_07404_),
    .A1(_07405_),
    .A2(_07406_),
    .A3(_07407_),
    .S0(net399),
    .S1(net397),
    .X(_07408_));
 sky130_fd_sc_hd__mux4_2 _19071_ (.A0(\w[33][20] ),
    .A1(\w[37][20] ),
    .A2(\w[35][20] ),
    .A3(\w[39][20] ),
    .S0(net538),
    .S1(net412),
    .X(_07409_));
 sky130_fd_sc_hd__mux4_2 _19072_ (.A0(\w[41][20] ),
    .A1(\w[45][20] ),
    .A2(\w[43][20] ),
    .A3(\w[47][20] ),
    .S0(net538),
    .S1(net412),
    .X(_07410_));
 sky130_fd_sc_hd__mux4_2 _19073_ (.A0(\w[49][20] ),
    .A1(\w[53][20] ),
    .A2(\w[51][20] ),
    .A3(\w[55][20] ),
    .S0(net538),
    .S1(net412),
    .X(_07411_));
 sky130_fd_sc_hd__mux4_2 _19074_ (.A0(\w[57][20] ),
    .A1(\w[61][20] ),
    .A2(\w[59][20] ),
    .A3(\w[63][20] ),
    .S0(net538),
    .S1(net412),
    .X(_07412_));
 sky130_fd_sc_hd__mux4_2 _19075_ (.A0(_07409_),
    .A1(_07410_),
    .A2(_07411_),
    .A3(_07412_),
    .S0(net399),
    .S1(net397),
    .X(_07413_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1057 ();
 sky130_fd_sc_hd__mux2i_4 _19077_ (.A0(_07408_),
    .A1(_07413_),
    .S(\count7_1[5] ),
    .Y(_11740_));
 sky130_fd_sc_hd__mux4_2 _19078_ (.A0(\w[1][21] ),
    .A1(\w[5][21] ),
    .A2(\w[3][21] ),
    .A3(\w[7][21] ),
    .S0(net403),
    .S1(net411),
    .X(_07415_));
 sky130_fd_sc_hd__mux4_2 _19079_ (.A0(\w[9][21] ),
    .A1(\w[13][21] ),
    .A2(\w[11][21] ),
    .A3(\w[15][21] ),
    .S0(net403),
    .S1(net411),
    .X(_07416_));
 sky130_fd_sc_hd__mux4_2 _19080_ (.A0(\w[17][21] ),
    .A1(\w[21][21] ),
    .A2(\w[19][21] ),
    .A3(\w[23][21] ),
    .S0(net402),
    .S1(net410),
    .X(_07417_));
 sky130_fd_sc_hd__mux4_2 _19081_ (.A0(\w[25][21] ),
    .A1(\w[29][21] ),
    .A2(\w[27][21] ),
    .A3(\w[31][21] ),
    .S0(net402),
    .S1(net410),
    .X(_07418_));
 sky130_fd_sc_hd__mux4_2 _19082_ (.A0(_07415_),
    .A1(_07416_),
    .A2(_07417_),
    .A3(_07418_),
    .S0(net399),
    .S1(net397),
    .X(_07419_));
 sky130_fd_sc_hd__mux4_2 _19083_ (.A0(\w[33][21] ),
    .A1(\w[37][21] ),
    .A2(\w[35][21] ),
    .A3(\w[39][21] ),
    .S0(net402),
    .S1(net410),
    .X(_07420_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1056 ();
 sky130_fd_sc_hd__mux4_2 _19085_ (.A0(\w[41][21] ),
    .A1(\w[45][21] ),
    .A2(\w[43][21] ),
    .A3(\w[47][21] ),
    .S0(net402),
    .S1(net410),
    .X(_07422_));
 sky130_fd_sc_hd__mux4_2 _19086_ (.A0(\w[49][21] ),
    .A1(\w[53][21] ),
    .A2(\w[51][21] ),
    .A3(\w[55][21] ),
    .S0(net402),
    .S1(net410),
    .X(_07423_));
 sky130_fd_sc_hd__mux4_2 _19087_ (.A0(\w[57][21] ),
    .A1(\w[61][21] ),
    .A2(\w[59][21] ),
    .A3(\w[63][21] ),
    .S0(net402),
    .S1(net410),
    .X(_07424_));
 sky130_fd_sc_hd__mux4_2 _19088_ (.A0(_07420_),
    .A1(_07422_),
    .A2(_07423_),
    .A3(_07424_),
    .S0(net399),
    .S1(net397),
    .X(_07425_));
 sky130_fd_sc_hd__mux2i_4 _19089_ (.A0(_07419_),
    .A1(_07425_),
    .S(net394),
    .Y(_11748_));
 sky130_fd_sc_hd__mux4_2 _19090_ (.A0(\w[1][22] ),
    .A1(\w[5][22] ),
    .A2(\w[3][22] ),
    .A3(\w[7][22] ),
    .S0(net403),
    .S1(net411),
    .X(_07426_));
 sky130_fd_sc_hd__mux4_2 _19091_ (.A0(\w[9][22] ),
    .A1(\w[13][22] ),
    .A2(\w[11][22] ),
    .A3(\w[15][22] ),
    .S0(net403),
    .S1(net411),
    .X(_07427_));
 sky130_fd_sc_hd__mux4_2 _19092_ (.A0(\w[17][22] ),
    .A1(\w[21][22] ),
    .A2(\w[19][22] ),
    .A3(\w[23][22] ),
    .S0(net403),
    .S1(net411),
    .X(_07428_));
 sky130_fd_sc_hd__mux4_2 _19093_ (.A0(\w[25][22] ),
    .A1(\w[29][22] ),
    .A2(\w[27][22] ),
    .A3(\w[31][22] ),
    .S0(net403),
    .S1(net411),
    .X(_07429_));
 sky130_fd_sc_hd__mux4_2 _19094_ (.A0(_07426_),
    .A1(_07427_),
    .A2(_07428_),
    .A3(_07429_),
    .S0(net399),
    .S1(net397),
    .X(_07430_));
 sky130_fd_sc_hd__mux4_2 _19095_ (.A0(\w[33][22] ),
    .A1(\w[37][22] ),
    .A2(\w[35][22] ),
    .A3(\w[39][22] ),
    .S0(net403),
    .S1(net411),
    .X(_07431_));
 sky130_fd_sc_hd__mux4_2 _19096_ (.A0(\w[41][22] ),
    .A1(\w[45][22] ),
    .A2(\w[43][22] ),
    .A3(\w[47][22] ),
    .S0(net403),
    .S1(net411),
    .X(_07432_));
 sky130_fd_sc_hd__mux4_2 _19097_ (.A0(\w[49][22] ),
    .A1(\w[53][22] ),
    .A2(\w[51][22] ),
    .A3(\w[55][22] ),
    .S0(net403),
    .S1(net411),
    .X(_07433_));
 sky130_fd_sc_hd__mux4_2 _19098_ (.A0(\w[57][22] ),
    .A1(\w[61][22] ),
    .A2(\w[59][22] ),
    .A3(\w[63][22] ),
    .S0(net403),
    .S1(net411),
    .X(_07434_));
 sky130_fd_sc_hd__mux4_2 _19099_ (.A0(_07431_),
    .A1(_07432_),
    .A2(_07433_),
    .A3(_07434_),
    .S0(net399),
    .S1(net397),
    .X(_07435_));
 sky130_fd_sc_hd__mux2i_4 _19100_ (.A0(_07430_),
    .A1(_07435_),
    .S(net394),
    .Y(_11756_));
 sky130_fd_sc_hd__mux4_2 _19101_ (.A0(\w[1][23] ),
    .A1(\w[5][23] ),
    .A2(\w[3][23] ),
    .A3(\w[7][23] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07436_));
 sky130_fd_sc_hd__mux4_2 _19102_ (.A0(\w[9][23] ),
    .A1(\w[13][23] ),
    .A2(\w[11][23] ),
    .A3(\w[15][23] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07437_));
 sky130_fd_sc_hd__mux4_2 _19103_ (.A0(\w[17][23] ),
    .A1(\w[21][23] ),
    .A2(\w[19][23] ),
    .A3(\w[23][23] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07438_));
 sky130_fd_sc_hd__mux4_2 _19104_ (.A0(\w[25][23] ),
    .A1(\w[29][23] ),
    .A2(\w[27][23] ),
    .A3(\w[31][23] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07439_));
 sky130_fd_sc_hd__mux4_2 _19105_ (.A0(_07436_),
    .A1(_07437_),
    .A2(_07438_),
    .A3(_07439_),
    .S0(net400),
    .S1(\count7_1[4] ),
    .X(_07440_));
 sky130_fd_sc_hd__mux4_2 _19106_ (.A0(\w[33][23] ),
    .A1(\w[37][23] ),
    .A2(\w[35][23] ),
    .A3(\w[39][23] ),
    .S0(net406),
    .S1(net412),
    .X(_07441_));
 sky130_fd_sc_hd__mux4_2 _19107_ (.A0(\w[41][23] ),
    .A1(\w[45][23] ),
    .A2(\w[43][23] ),
    .A3(\w[47][23] ),
    .S0(net406),
    .S1(net412),
    .X(_07442_));
 sky130_fd_sc_hd__mux4_2 _19108_ (.A0(\w[49][23] ),
    .A1(\w[53][23] ),
    .A2(\w[51][23] ),
    .A3(\w[55][23] ),
    .S0(net406),
    .S1(net412),
    .X(_07443_));
 sky130_fd_sc_hd__mux4_2 _19109_ (.A0(\w[57][23] ),
    .A1(\w[61][23] ),
    .A2(\w[59][23] ),
    .A3(\w[63][23] ),
    .S0(net406),
    .S1(net412),
    .X(_07444_));
 sky130_fd_sc_hd__mux4_2 _19110_ (.A0(_07441_),
    .A1(_07442_),
    .A2(_07443_),
    .A3(_07444_),
    .S0(net537),
    .S1(net396),
    .X(_07445_));
 sky130_fd_sc_hd__mux2i_4 _19111_ (.A0(_07440_),
    .A1(_07445_),
    .S(net395),
    .Y(_11764_));
 sky130_fd_sc_hd__mux4_2 _19112_ (.A0(\w[1][24] ),
    .A1(\w[5][24] ),
    .A2(\w[3][24] ),
    .A3(\w[7][24] ),
    .S0(net401),
    .S1(net408),
    .X(_07446_));
 sky130_fd_sc_hd__mux4_2 _19113_ (.A0(\w[9][24] ),
    .A1(\w[13][24] ),
    .A2(\w[11][24] ),
    .A3(\w[15][24] ),
    .S0(net401),
    .S1(net408),
    .X(_07447_));
 sky130_fd_sc_hd__mux4_2 _19114_ (.A0(\w[17][24] ),
    .A1(\w[21][24] ),
    .A2(\w[19][24] ),
    .A3(\w[23][24] ),
    .S0(net401),
    .S1(net408),
    .X(_07448_));
 sky130_fd_sc_hd__mux4_2 _19115_ (.A0(\w[25][24] ),
    .A1(\w[29][24] ),
    .A2(\w[27][24] ),
    .A3(\w[31][24] ),
    .S0(net401),
    .S1(net408),
    .X(_07449_));
 sky130_fd_sc_hd__mux4_2 _19116_ (.A0(_07446_),
    .A1(_07447_),
    .A2(_07448_),
    .A3(_07449_),
    .S0(net398),
    .S1(net396),
    .X(_07450_));
 sky130_fd_sc_hd__mux4_2 _19117_ (.A0(\w[33][24] ),
    .A1(\w[37][24] ),
    .A2(\w[35][24] ),
    .A3(\w[39][24] ),
    .S0(net404),
    .S1(net411),
    .X(_07451_));
 sky130_fd_sc_hd__mux4_2 _19118_ (.A0(\w[41][24] ),
    .A1(\w[45][24] ),
    .A2(\w[43][24] ),
    .A3(\w[47][24] ),
    .S0(net404),
    .S1(net411),
    .X(_07452_));
 sky130_fd_sc_hd__mux4_2 _19119_ (.A0(\w[49][24] ),
    .A1(\w[53][24] ),
    .A2(\w[51][24] ),
    .A3(\w[55][24] ),
    .S0(net404),
    .S1(net411),
    .X(_07453_));
 sky130_fd_sc_hd__mux4_2 _19120_ (.A0(\w[57][24] ),
    .A1(\w[61][24] ),
    .A2(\w[59][24] ),
    .A3(\w[63][24] ),
    .S0(net404),
    .S1(net410),
    .X(_07454_));
 sky130_fd_sc_hd__mux4_2 _19121_ (.A0(_07451_),
    .A1(_07452_),
    .A2(_07453_),
    .A3(_07454_),
    .S0(net537),
    .S1(net396),
    .X(_07455_));
 sky130_fd_sc_hd__mux2i_4 _19122_ (.A0(_07450_),
    .A1(_07455_),
    .S(net394),
    .Y(_11772_));
 sky130_fd_sc_hd__mux4_2 _19123_ (.A0(\w[1][25] ),
    .A1(\w[5][25] ),
    .A2(\w[3][25] ),
    .A3(\w[7][25] ),
    .S0(net403),
    .S1(net411),
    .X(_07456_));
 sky130_fd_sc_hd__mux4_2 _19124_ (.A0(\w[9][25] ),
    .A1(\w[13][25] ),
    .A2(\w[11][25] ),
    .A3(\w[15][25] ),
    .S0(net403),
    .S1(net411),
    .X(_07457_));
 sky130_fd_sc_hd__mux4_2 _19125_ (.A0(\w[17][25] ),
    .A1(\w[21][25] ),
    .A2(\w[19][25] ),
    .A3(\w[23][25] ),
    .S0(net403),
    .S1(net411),
    .X(_07458_));
 sky130_fd_sc_hd__mux4_2 _19126_ (.A0(\w[25][25] ),
    .A1(\w[29][25] ),
    .A2(\w[27][25] ),
    .A3(\w[31][25] ),
    .S0(net403),
    .S1(net411),
    .X(_07459_));
 sky130_fd_sc_hd__mux4_2 _19127_ (.A0(_07456_),
    .A1(_07457_),
    .A2(_07458_),
    .A3(_07459_),
    .S0(net398),
    .S1(net397),
    .X(_07460_));
 sky130_fd_sc_hd__mux4_2 _19128_ (.A0(\w[33][25] ),
    .A1(\w[37][25] ),
    .A2(\w[35][25] ),
    .A3(\w[39][25] ),
    .S0(net403),
    .S1(net411),
    .X(_07461_));
 sky130_fd_sc_hd__mux4_2 _19129_ (.A0(\w[41][25] ),
    .A1(\w[45][25] ),
    .A2(\w[43][25] ),
    .A3(\w[47][25] ),
    .S0(net403),
    .S1(net411),
    .X(_07462_));
 sky130_fd_sc_hd__mux4_2 _19130_ (.A0(\w[49][25] ),
    .A1(\w[53][25] ),
    .A2(\w[51][25] ),
    .A3(\w[55][25] ),
    .S0(net403),
    .S1(net411),
    .X(_07463_));
 sky130_fd_sc_hd__mux4_2 _19131_ (.A0(\w[57][25] ),
    .A1(\w[61][25] ),
    .A2(\w[59][25] ),
    .A3(\w[63][25] ),
    .S0(net403),
    .S1(net411),
    .X(_07464_));
 sky130_fd_sc_hd__mux4_2 _19132_ (.A0(_07461_),
    .A1(_07462_),
    .A2(_07463_),
    .A3(_07464_),
    .S0(net537),
    .S1(net397),
    .X(_07465_));
 sky130_fd_sc_hd__mux2i_4 _19133_ (.A0(_07460_),
    .A1(_07465_),
    .S(net394),
    .Y(_11780_));
 sky130_fd_sc_hd__mux4_2 _19134_ (.A0(\w[1][26] ),
    .A1(\w[5][26] ),
    .A2(\w[3][26] ),
    .A3(\w[7][26] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07466_));
 sky130_fd_sc_hd__mux4_2 _19135_ (.A0(\w[9][26] ),
    .A1(\w[13][26] ),
    .A2(\w[11][26] ),
    .A3(\w[15][26] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07467_));
 sky130_fd_sc_hd__mux4_2 _19136_ (.A0(\w[17][26] ),
    .A1(\w[21][26] ),
    .A2(\w[19][26] ),
    .A3(\w[23][26] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07468_));
 sky130_fd_sc_hd__mux4_2 _19137_ (.A0(\w[25][26] ),
    .A1(\w[29][26] ),
    .A2(\w[27][26] ),
    .A3(\w[31][26] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07469_));
 sky130_fd_sc_hd__mux4_2 _19138_ (.A0(_07466_),
    .A1(_07467_),
    .A2(_07468_),
    .A3(_07469_),
    .S0(net400),
    .S1(\count7_1[4] ),
    .X(_07470_));
 sky130_fd_sc_hd__mux4_2 _19139_ (.A0(\w[33][26] ),
    .A1(\w[37][26] ),
    .A2(\w[35][26] ),
    .A3(\w[39][26] ),
    .S0(net405),
    .S1(net409),
    .X(_07471_));
 sky130_fd_sc_hd__mux4_2 _19140_ (.A0(\w[41][26] ),
    .A1(\w[45][26] ),
    .A2(\w[43][26] ),
    .A3(\w[47][26] ),
    .S0(net405),
    .S1(net409),
    .X(_07472_));
 sky130_fd_sc_hd__mux4_2 _19141_ (.A0(\w[49][26] ),
    .A1(\w[53][26] ),
    .A2(\w[51][26] ),
    .A3(\w[55][26] ),
    .S0(net405),
    .S1(net409),
    .X(_07473_));
 sky130_fd_sc_hd__mux4_2 _19142_ (.A0(\w[57][26] ),
    .A1(\w[61][26] ),
    .A2(\w[59][26] ),
    .A3(\w[63][26] ),
    .S0(net405),
    .S1(net409),
    .X(_07474_));
 sky130_fd_sc_hd__mux4_2 _19143_ (.A0(_07471_),
    .A1(_07472_),
    .A2(_07473_),
    .A3(_07474_),
    .S0(net400),
    .S1(net536),
    .X(_07475_));
 sky130_fd_sc_hd__mux2i_4 _19144_ (.A0(_07470_),
    .A1(_07475_),
    .S(net395),
    .Y(_11788_));
 sky130_fd_sc_hd__mux4_2 _19145_ (.A0(\w[1][27] ),
    .A1(\w[5][27] ),
    .A2(\w[3][27] ),
    .A3(\w[7][27] ),
    .S0(net401),
    .S1(net408),
    .X(_07476_));
 sky130_fd_sc_hd__mux4_2 _19146_ (.A0(\w[9][27] ),
    .A1(\w[13][27] ),
    .A2(\w[11][27] ),
    .A3(\w[15][27] ),
    .S0(net401),
    .S1(net408),
    .X(_07477_));
 sky130_fd_sc_hd__mux4_2 _19147_ (.A0(\w[17][27] ),
    .A1(\w[21][27] ),
    .A2(\w[19][27] ),
    .A3(\w[23][27] ),
    .S0(net401),
    .S1(net408),
    .X(_07478_));
 sky130_fd_sc_hd__mux4_2 _19148_ (.A0(\w[25][27] ),
    .A1(\w[29][27] ),
    .A2(\w[27][27] ),
    .A3(\w[31][27] ),
    .S0(net401),
    .S1(net408),
    .X(_07479_));
 sky130_fd_sc_hd__mux4_2 _19149_ (.A0(_07476_),
    .A1(_07477_),
    .A2(_07478_),
    .A3(_07479_),
    .S0(net398),
    .S1(net396),
    .X(_07480_));
 sky130_fd_sc_hd__mux4_2 _19150_ (.A0(\w[33][27] ),
    .A1(\w[37][27] ),
    .A2(\w[35][27] ),
    .A3(\w[39][27] ),
    .S0(net406),
    .S1(net412),
    .X(_07481_));
 sky130_fd_sc_hd__mux4_2 _19151_ (.A0(\w[41][27] ),
    .A1(\w[45][27] ),
    .A2(\w[43][27] ),
    .A3(\w[47][27] ),
    .S0(net406),
    .S1(net412),
    .X(_07482_));
 sky130_fd_sc_hd__mux4_2 _19152_ (.A0(\w[49][27] ),
    .A1(\w[53][27] ),
    .A2(\w[51][27] ),
    .A3(\w[55][27] ),
    .S0(net406),
    .S1(net412),
    .X(_07483_));
 sky130_fd_sc_hd__mux4_2 _19153_ (.A0(\w[57][27] ),
    .A1(\w[61][27] ),
    .A2(\w[59][27] ),
    .A3(\w[63][27] ),
    .S0(net406),
    .S1(net412),
    .X(_07484_));
 sky130_fd_sc_hd__mux4_2 _19154_ (.A0(_07481_),
    .A1(_07482_),
    .A2(_07483_),
    .A3(_07484_),
    .S0(net398),
    .S1(net396),
    .X(_07485_));
 sky130_fd_sc_hd__mux2i_4 _19155_ (.A0(_07480_),
    .A1(_07485_),
    .S(net394),
    .Y(_11796_));
 sky130_fd_sc_hd__mux4_2 _19156_ (.A0(\w[1][28] ),
    .A1(\w[5][28] ),
    .A2(\w[3][28] ),
    .A3(\w[7][28] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07486_));
 sky130_fd_sc_hd__mux4_2 _19157_ (.A0(\w[9][28] ),
    .A1(\w[13][28] ),
    .A2(\w[11][28] ),
    .A3(\w[15][28] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07487_));
 sky130_fd_sc_hd__mux4_2 _19158_ (.A0(\w[17][28] ),
    .A1(\w[21][28] ),
    .A2(\w[19][28] ),
    .A3(\w[23][28] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07488_));
 sky130_fd_sc_hd__mux4_2 _19159_ (.A0(\w[25][28] ),
    .A1(\w[29][28] ),
    .A2(\w[27][28] ),
    .A3(\w[31][28] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07489_));
 sky130_fd_sc_hd__mux4_2 _19160_ (.A0(_07486_),
    .A1(_07487_),
    .A2(_07488_),
    .A3(_07489_),
    .S0(net400),
    .S1(\count7_1[4] ),
    .X(_07490_));
 sky130_fd_sc_hd__mux4_2 _19161_ (.A0(\w[33][28] ),
    .A1(\w[37][28] ),
    .A2(\w[35][28] ),
    .A3(\w[39][28] ),
    .S0(net407),
    .S1(net409),
    .X(_07491_));
 sky130_fd_sc_hd__mux4_2 _19162_ (.A0(\w[41][28] ),
    .A1(\w[45][28] ),
    .A2(\w[43][28] ),
    .A3(\w[47][28] ),
    .S0(net407),
    .S1(net409),
    .X(_07492_));
 sky130_fd_sc_hd__mux4_2 _19163_ (.A0(\w[49][28] ),
    .A1(\w[53][28] ),
    .A2(\w[51][28] ),
    .A3(\w[55][28] ),
    .S0(net407),
    .S1(net409),
    .X(_07493_));
 sky130_fd_sc_hd__mux4_2 _19164_ (.A0(\w[57][28] ),
    .A1(\w[61][28] ),
    .A2(\w[59][28] ),
    .A3(\w[63][28] ),
    .S0(net407),
    .S1(net409),
    .X(_07494_));
 sky130_fd_sc_hd__mux4_2 _19165_ (.A0(_07491_),
    .A1(_07492_),
    .A2(_07493_),
    .A3(_07494_),
    .S0(net400),
    .S1(net536),
    .X(_07495_));
 sky130_fd_sc_hd__mux2i_4 _19166_ (.A0(_07490_),
    .A1(_07495_),
    .S(net395),
    .Y(_11804_));
 sky130_fd_sc_hd__mux4_2 _19167_ (.A0(\w[1][29] ),
    .A1(\w[5][29] ),
    .A2(\w[3][29] ),
    .A3(\w[7][29] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07496_));
 sky130_fd_sc_hd__mux4_2 _19168_ (.A0(\w[9][29] ),
    .A1(\w[13][29] ),
    .A2(\w[11][29] ),
    .A3(\w[15][29] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07497_));
 sky130_fd_sc_hd__mux4_2 _19169_ (.A0(\w[17][29] ),
    .A1(\w[21][29] ),
    .A2(\w[19][29] ),
    .A3(\w[23][29] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07498_));
 sky130_fd_sc_hd__mux4_2 _19170_ (.A0(\w[25][29] ),
    .A1(\w[29][29] ),
    .A2(\w[27][29] ),
    .A3(\w[31][29] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07499_));
 sky130_fd_sc_hd__mux4_2 _19171_ (.A0(_07496_),
    .A1(_07497_),
    .A2(_07498_),
    .A3(_07499_),
    .S0(net400),
    .S1(\count7_1[4] ),
    .X(_07500_));
 sky130_fd_sc_hd__mux4_2 _19172_ (.A0(\w[33][29] ),
    .A1(\w[37][29] ),
    .A2(\w[35][29] ),
    .A3(\w[39][29] ),
    .S0(net406),
    .S1(net412),
    .X(_07501_));
 sky130_fd_sc_hd__mux4_2 _19173_ (.A0(\w[41][29] ),
    .A1(\w[45][29] ),
    .A2(\w[43][29] ),
    .A3(\w[47][29] ),
    .S0(net406),
    .S1(net412),
    .X(_07502_));
 sky130_fd_sc_hd__mux4_2 _19174_ (.A0(\w[49][29] ),
    .A1(\w[53][29] ),
    .A2(\w[51][29] ),
    .A3(\w[55][29] ),
    .S0(net406),
    .S1(net412),
    .X(_07503_));
 sky130_fd_sc_hd__mux4_2 _19175_ (.A0(\w[57][29] ),
    .A1(\w[61][29] ),
    .A2(\w[59][29] ),
    .A3(\w[63][29] ),
    .S0(net406),
    .S1(net412),
    .X(_07504_));
 sky130_fd_sc_hd__mux4_2 _19176_ (.A0(_07501_),
    .A1(_07502_),
    .A2(_07503_),
    .A3(_07504_),
    .S0(net537),
    .S1(net536),
    .X(_07505_));
 sky130_fd_sc_hd__mux2i_4 _19177_ (.A0(_07500_),
    .A1(_07505_),
    .S(\count7_1[5] ),
    .Y(_11812_));
 sky130_fd_sc_hd__mux4_2 _19178_ (.A0(\w[1][30] ),
    .A1(\w[5][30] ),
    .A2(\w[3][30] ),
    .A3(\w[7][30] ),
    .S0(net407),
    .S1(net409),
    .X(_07506_));
 sky130_fd_sc_hd__mux4_2 _19179_ (.A0(\w[9][30] ),
    .A1(\w[13][30] ),
    .A2(\w[11][30] ),
    .A3(\w[15][30] ),
    .S0(net407),
    .S1(net409),
    .X(_07507_));
 sky130_fd_sc_hd__mux4_2 _19180_ (.A0(\w[17][30] ),
    .A1(\w[21][30] ),
    .A2(\w[19][30] ),
    .A3(\w[23][30] ),
    .S0(net407),
    .S1(\count7_1[1] ),
    .X(_07508_));
 sky130_fd_sc_hd__mux4_2 _19181_ (.A0(\w[25][30] ),
    .A1(\w[29][30] ),
    .A2(\w[27][30] ),
    .A3(\w[31][30] ),
    .S0(net407),
    .S1(net409),
    .X(_07509_));
 sky130_fd_sc_hd__mux4_2 _19182_ (.A0(_07506_),
    .A1(_07507_),
    .A2(_07508_),
    .A3(_07509_),
    .S0(net400),
    .S1(\count7_1[4] ),
    .X(_07510_));
 sky130_fd_sc_hd__mux4_2 _19183_ (.A0(\w[33][30] ),
    .A1(\w[37][30] ),
    .A2(\w[35][30] ),
    .A3(\w[39][30] ),
    .S0(net538),
    .S1(net412),
    .X(_07511_));
 sky130_fd_sc_hd__mux4_2 _19184_ (.A0(\w[41][30] ),
    .A1(\w[45][30] ),
    .A2(\w[43][30] ),
    .A3(\w[47][30] ),
    .S0(net538),
    .S1(net412),
    .X(_07512_));
 sky130_fd_sc_hd__mux4_2 _19185_ (.A0(\w[49][30] ),
    .A1(\w[53][30] ),
    .A2(\w[51][30] ),
    .A3(\w[55][30] ),
    .S0(net538),
    .S1(net412),
    .X(_07513_));
 sky130_fd_sc_hd__mux4_2 _19186_ (.A0(\w[57][30] ),
    .A1(\w[61][30] ),
    .A2(\w[59][30] ),
    .A3(\w[63][30] ),
    .S0(net538),
    .S1(net412),
    .X(_07514_));
 sky130_fd_sc_hd__mux4_2 _19187_ (.A0(_07511_),
    .A1(_07512_),
    .A2(_07513_),
    .A3(_07514_),
    .S0(net399),
    .S1(net397),
    .X(_07515_));
 sky130_fd_sc_hd__mux2i_2 _19188_ (.A0(_07510_),
    .A1(_07515_),
    .S(\count7_1[5] ),
    .Y(_11820_));
 sky130_fd_sc_hd__inv_1 _19189_ (.A(\hash.CA1.w_i2[1] ),
    .Y(_12367_));
 sky130_fd_sc_hd__clkinv_1 _19190_ (.A(\hash.CA1.w_i2[0] ),
    .Y(_12372_));
 sky130_fd_sc_hd__inv_1 _19191_ (.A(\hash.CA1.w_i2[3] ),
    .Y(_12382_));
 sky130_fd_sc_hd__inv_2 _19192_ (.A(\hash.CA1.w_i2[5] ),
    .Y(_12390_));
 sky130_fd_sc_hd__inv_1 _19193_ (.A(\hash.CA1.w_i2[7] ),
    .Y(_12398_));
 sky130_fd_sc_hd__clkinv_2 _19194_ (.A(\hash.CA1.w_i2[8] ),
    .Y(_12403_));
 sky130_fd_sc_hd__inv_1 _19195_ (.A(\hash.CA1.w_i2[11] ),
    .Y(_12414_));
 sky130_fd_sc_hd__inv_1 _19196_ (.A(\hash.CA1.w_i2[12] ),
    .Y(_12419_));
 sky130_fd_sc_hd__inv_4 _19197_ (.A(\hash.CA1.w_i2[14] ),
    .Y(_12427_));
 sky130_fd_sc_hd__inv_4 _19198_ (.A(\hash.CA1.w_i2[15] ),
    .Y(_12432_));
 sky130_fd_sc_hd__inv_4 _19199_ (.A(\hash.CA1.w_i2[16] ),
    .Y(_12437_));
 sky130_fd_sc_hd__inv_1 _19200_ (.A(\hash.CA1.w_i2[17] ),
    .Y(_12442_));
 sky130_fd_sc_hd__clkinvlp_2 _19201_ (.A(\hash.CA1.w_i2[23] ),
    .Y(_12462_));
 sky130_fd_sc_hd__inv_4 _19202_ (.A(\hash.CA1.w_i2[24] ),
    .Y(_12467_));
 sky130_fd_sc_hd__inv_4 _19203_ (.A(\hash.CA1.w_i2[25] ),
    .Y(_12472_));
 sky130_fd_sc_hd__inv_1 _19204_ (.A(\hash.CA1.w_i2[26] ),
    .Y(_12477_));
 sky130_fd_sc_hd__inv_6 _19205_ (.A(\hash.CA1.w_i2[27] ),
    .Y(_12482_));
 sky130_fd_sc_hd__inv_1 _19206_ (.A(\hash.CA1.w_i2[28] ),
    .Y(_12487_));
 sky130_fd_sc_hd__inv_1 _19207_ (.A(_12725_),
    .Y(_12727_));
 sky130_fd_sc_hd__clkinv_2 _19208_ (.A(_06771_),
    .Y(_12793_));
 sky130_fd_sc_hd__inv_1 _19209_ (.A(_12898_),
    .Y(_12894_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1052 ();
 sky130_fd_sc_hd__mux4_2 _19214_ (.A0(\w[0][0] ),
    .A1(\w[4][0] ),
    .A2(\w[2][0] ),
    .A3(\w[6][0] ),
    .S0(net479),
    .S1(net489),
    .X(_07520_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1048 ();
 sky130_fd_sc_hd__mux4_2 _19219_ (.A0(\w[8][0] ),
    .A1(\w[12][0] ),
    .A2(\w[10][0] ),
    .A3(\w[14][0] ),
    .S0(net479),
    .S1(net489),
    .X(_07525_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1046 ();
 sky130_fd_sc_hd__mux4_2 _19222_ (.A0(\w[16][0] ),
    .A1(\w[20][0] ),
    .A2(\w[18][0] ),
    .A3(\w[22][0] ),
    .S0(net479),
    .S1(net489),
    .X(_07528_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1043 ();
 sky130_fd_sc_hd__mux4_2 _19226_ (.A0(\w[24][0] ),
    .A1(\w[28][0] ),
    .A2(\w[26][0] ),
    .A3(\w[30][0] ),
    .S0(net479),
    .S1(net489),
    .X(_07532_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1039 ();
 sky130_fd_sc_hd__mux4_2 _19231_ (.A0(_07520_),
    .A1(_07525_),
    .A2(_07528_),
    .A3(_07532_),
    .S0(net477),
    .S1(net475),
    .X(_07537_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1037 ();
 sky130_fd_sc_hd__mux4_2 _19234_ (.A0(\w[32][0] ),
    .A1(\w[36][0] ),
    .A2(\w[34][0] ),
    .A3(\w[38][0] ),
    .S0(net484),
    .S1(net490),
    .X(_07540_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1035 ();
 sky130_fd_sc_hd__mux4_2 _19237_ (.A0(\w[40][0] ),
    .A1(\w[44][0] ),
    .A2(\w[42][0] ),
    .A3(\w[46][0] ),
    .S0(net484),
    .S1(net490),
    .X(_07543_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1033 ();
 sky130_fd_sc_hd__mux4_2 _19240_ (.A0(\w[48][0] ),
    .A1(\w[52][0] ),
    .A2(\w[50][0] ),
    .A3(\w[54][0] ),
    .S0(net484),
    .S1(net490),
    .X(_07546_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1031 ();
 sky130_fd_sc_hd__mux4_2 _19243_ (.A0(\w[56][0] ),
    .A1(\w[60][0] ),
    .A2(\w[58][0] ),
    .A3(\w[62][0] ),
    .S0(net484),
    .S1(net490),
    .X(_07549_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1029 ();
 sky130_fd_sc_hd__mux4_2 _19246_ (.A0(_07540_),
    .A1(_07543_),
    .A2(_07546_),
    .A3(_07549_),
    .S0(net477),
    .S1(net475),
    .X(_07552_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1028 ();
 sky130_fd_sc_hd__mux2i_4 _19248_ (.A0(_07537_),
    .A1(_07552_),
    .S(net472),
    .Y(_11581_));
 sky130_fd_sc_hd__mux4_2 _19249_ (.A0(\w[0][1] ),
    .A1(\w[4][1] ),
    .A2(\w[2][1] ),
    .A3(\w[6][1] ),
    .S0(net479),
    .S1(net489),
    .X(_07554_));
 sky130_fd_sc_hd__mux4_2 _19250_ (.A0(\w[8][1] ),
    .A1(\w[12][1] ),
    .A2(\w[10][1] ),
    .A3(\w[14][1] ),
    .S0(net479),
    .S1(net489),
    .X(_07555_));
 sky130_fd_sc_hd__mux4_2 _19251_ (.A0(\w[16][1] ),
    .A1(\w[20][1] ),
    .A2(\w[18][1] ),
    .A3(\w[22][1] ),
    .S0(net479),
    .S1(net489),
    .X(_07556_));
 sky130_fd_sc_hd__mux4_2 _19252_ (.A0(\w[24][1] ),
    .A1(\w[28][1] ),
    .A2(\w[26][1] ),
    .A3(\w[30][1] ),
    .S0(net479),
    .S1(net489),
    .X(_07557_));
 sky130_fd_sc_hd__mux4_2 _19253_ (.A0(_07554_),
    .A1(_07555_),
    .A2(_07556_),
    .A3(_07557_),
    .S0(net477),
    .S1(net475),
    .X(_07558_));
 sky130_fd_sc_hd__mux4_2 _19254_ (.A0(\w[32][1] ),
    .A1(\w[36][1] ),
    .A2(\w[34][1] ),
    .A3(\w[38][1] ),
    .S0(net484),
    .S1(net490),
    .X(_07559_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1027 ();
 sky130_fd_sc_hd__mux4_2 _19256_ (.A0(\w[40][1] ),
    .A1(\w[44][1] ),
    .A2(\w[42][1] ),
    .A3(\w[46][1] ),
    .S0(net484),
    .S1(net490),
    .X(_07561_));
 sky130_fd_sc_hd__mux4_2 _19257_ (.A0(\w[48][1] ),
    .A1(\w[52][1] ),
    .A2(\w[50][1] ),
    .A3(\w[54][1] ),
    .S0(net484),
    .S1(net490),
    .X(_07562_));
 sky130_fd_sc_hd__mux4_2 _19258_ (.A0(\w[56][1] ),
    .A1(\w[60][1] ),
    .A2(\w[58][1] ),
    .A3(\w[62][1] ),
    .S0(net484),
    .S1(net490),
    .X(_07563_));
 sky130_fd_sc_hd__mux4_2 _19259_ (.A0(_07559_),
    .A1(_07561_),
    .A2(_07562_),
    .A3(_07563_),
    .S0(net477),
    .S1(net475),
    .X(_07564_));
 sky130_fd_sc_hd__mux2i_4 _19260_ (.A0(_07558_),
    .A1(_07564_),
    .S(net472),
    .Y(_11586_));
 sky130_fd_sc_hd__mux4_2 _19261_ (.A0(\w[0][2] ),
    .A1(\w[4][2] ),
    .A2(\w[2][2] ),
    .A3(\w[6][2] ),
    .S0(net478),
    .S1(net486),
    .X(_07565_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1026 ();
 sky130_fd_sc_hd__mux4_2 _19263_ (.A0(\w[8][2] ),
    .A1(\w[12][2] ),
    .A2(\w[10][2] ),
    .A3(\w[14][2] ),
    .S0(net478),
    .S1(net486),
    .X(_07567_));
 sky130_fd_sc_hd__mux4_2 _19264_ (.A0(\w[16][2] ),
    .A1(\w[20][2] ),
    .A2(\w[18][2] ),
    .A3(\w[22][2] ),
    .S0(net478),
    .S1(net486),
    .X(_07568_));
 sky130_fd_sc_hd__mux4_2 _19265_ (.A0(\w[24][2] ),
    .A1(\w[28][2] ),
    .A2(\w[26][2] ),
    .A3(\w[30][2] ),
    .S0(net478),
    .S1(net486),
    .X(_07569_));
 sky130_fd_sc_hd__mux4_2 _19266_ (.A0(_07565_),
    .A1(_07567_),
    .A2(_07568_),
    .A3(_07569_),
    .S0(net476),
    .S1(net474),
    .X(_07570_));
 sky130_fd_sc_hd__mux4_2 _19267_ (.A0(\w[32][2] ),
    .A1(\w[36][2] ),
    .A2(\w[34][2] ),
    .A3(\w[38][2] ),
    .S0(net483),
    .S1(net491),
    .X(_07571_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1025 ();
 sky130_fd_sc_hd__mux4_2 _19269_ (.A0(\w[40][2] ),
    .A1(\w[44][2] ),
    .A2(\w[42][2] ),
    .A3(\w[46][2] ),
    .S0(net483),
    .S1(net491),
    .X(_07573_));
 sky130_fd_sc_hd__mux4_2 _19270_ (.A0(\w[48][2] ),
    .A1(\w[52][2] ),
    .A2(\w[50][2] ),
    .A3(\w[54][2] ),
    .S0(net483),
    .S1(net491),
    .X(_07574_));
 sky130_fd_sc_hd__mux4_2 _19271_ (.A0(\w[56][2] ),
    .A1(\w[60][2] ),
    .A2(\w[58][2] ),
    .A3(\w[62][2] ),
    .S0(net483),
    .S1(net491),
    .X(_07575_));
 sky130_fd_sc_hd__mux4_2 _19272_ (.A0(_07571_),
    .A1(_07573_),
    .A2(_07574_),
    .A3(_07575_),
    .S0(net546),
    .S1(net474),
    .X(_07576_));
 sky130_fd_sc_hd__mux2i_4 _19273_ (.A0(_07570_),
    .A1(_07576_),
    .S(net545),
    .Y(_11594_));
 sky130_fd_sc_hd__mux4_2 _19274_ (.A0(\w[0][3] ),
    .A1(\w[4][3] ),
    .A2(\w[2][3] ),
    .A3(\w[6][3] ),
    .S0(net485),
    .S1(\count16_1[1] ),
    .X(_07577_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1024 ();
 sky130_fd_sc_hd__mux4_2 _19276_ (.A0(\w[8][3] ),
    .A1(\w[12][3] ),
    .A2(\w[10][3] ),
    .A3(\w[14][3] ),
    .S0(net485),
    .S1(\count16_1[1] ),
    .X(_07579_));
 sky130_fd_sc_hd__mux4_2 _19277_ (.A0(\w[16][3] ),
    .A1(\w[20][3] ),
    .A2(\w[18][3] ),
    .A3(\w[22][3] ),
    .S0(net485),
    .S1(\count16_1[1] ),
    .X(_07580_));
 sky130_fd_sc_hd__mux4_2 _19278_ (.A0(\w[24][3] ),
    .A1(\w[28][3] ),
    .A2(\w[26][3] ),
    .A3(\w[30][3] ),
    .S0(net485),
    .S1(\count16_1[1] ),
    .X(_07581_));
 sky130_fd_sc_hd__mux4_2 _19279_ (.A0(_07577_),
    .A1(_07579_),
    .A2(_07580_),
    .A3(_07581_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07582_));
 sky130_fd_sc_hd__mux4_2 _19280_ (.A0(\w[32][3] ),
    .A1(\w[36][3] ),
    .A2(\w[34][3] ),
    .A3(\w[38][3] ),
    .S0(net485),
    .S1(net491),
    .X(_07583_));
 sky130_fd_sc_hd__mux4_2 _19281_ (.A0(\w[40][3] ),
    .A1(\w[44][3] ),
    .A2(\w[42][3] ),
    .A3(\w[46][3] ),
    .S0(net485),
    .S1(net491),
    .X(_07584_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1023 ();
 sky130_fd_sc_hd__mux4_2 _19283_ (.A0(\w[48][3] ),
    .A1(\w[52][3] ),
    .A2(\w[50][3] ),
    .A3(\w[54][3] ),
    .S0(net485),
    .S1(net491),
    .X(_07586_));
 sky130_fd_sc_hd__mux4_2 _19284_ (.A0(\w[56][3] ),
    .A1(\w[60][3] ),
    .A2(\w[58][3] ),
    .A3(\w[62][3] ),
    .S0(net485),
    .S1(net490),
    .X(_07587_));
 sky130_fd_sc_hd__mux4_2 _19285_ (.A0(_07583_),
    .A1(_07584_),
    .A2(_07586_),
    .A3(_07587_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07588_));
 sky130_fd_sc_hd__mux2i_4 _19286_ (.A0(_07582_),
    .A1(_07588_),
    .S(\count16_1[5] ),
    .Y(_11605_));
 sky130_fd_sc_hd__mux4_2 _19287_ (.A0(\w[0][4] ),
    .A1(\w[4][4] ),
    .A2(\w[2][4] ),
    .A3(\w[6][4] ),
    .S0(net478),
    .S1(net486),
    .X(_07589_));
 sky130_fd_sc_hd__mux4_2 _19288_ (.A0(\w[8][4] ),
    .A1(\w[12][4] ),
    .A2(\w[10][4] ),
    .A3(\w[14][4] ),
    .S0(net478),
    .S1(net486),
    .X(_07590_));
 sky130_fd_sc_hd__mux4_2 _19289_ (.A0(\w[16][4] ),
    .A1(\w[20][4] ),
    .A2(\w[18][4] ),
    .A3(\w[22][4] ),
    .S0(net478),
    .S1(net486),
    .X(_07591_));
 sky130_fd_sc_hd__mux4_2 _19290_ (.A0(\w[24][4] ),
    .A1(\w[28][4] ),
    .A2(\w[26][4] ),
    .A3(\w[30][4] ),
    .S0(net478),
    .S1(net486),
    .X(_07592_));
 sky130_fd_sc_hd__mux4_2 _19291_ (.A0(_07589_),
    .A1(_07590_),
    .A2(_07591_),
    .A3(_07592_),
    .S0(net546),
    .S1(net474),
    .X(_07593_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1022 ();
 sky130_fd_sc_hd__mux4_2 _19293_ (.A0(\w[32][4] ),
    .A1(\w[36][4] ),
    .A2(\w[34][4] ),
    .A3(\w[38][4] ),
    .S0(net478),
    .S1(net486),
    .X(_07595_));
 sky130_fd_sc_hd__mux4_2 _19294_ (.A0(\w[40][4] ),
    .A1(\w[44][4] ),
    .A2(\w[42][4] ),
    .A3(\w[46][4] ),
    .S0(net478),
    .S1(net486),
    .X(_07596_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1021 ();
 sky130_fd_sc_hd__mux4_2 _19296_ (.A0(\w[48][4] ),
    .A1(\w[52][4] ),
    .A2(\w[50][4] ),
    .A3(\w[54][4] ),
    .S0(net478),
    .S1(net486),
    .X(_07598_));
 sky130_fd_sc_hd__mux4_2 _19297_ (.A0(\w[56][4] ),
    .A1(\w[60][4] ),
    .A2(\w[58][4] ),
    .A3(\w[62][4] ),
    .S0(net478),
    .S1(net486),
    .X(_07599_));
 sky130_fd_sc_hd__mux4_2 _19298_ (.A0(_07595_),
    .A1(_07596_),
    .A2(_07598_),
    .A3(_07599_),
    .S0(net546),
    .S1(net474),
    .X(_07600_));
 sky130_fd_sc_hd__mux2i_4 _19299_ (.A0(_07593_),
    .A1(_07600_),
    .S(net545),
    .Y(_11613_));
 sky130_fd_sc_hd__mux4_2 _19300_ (.A0(\w[0][5] ),
    .A1(\w[4][5] ),
    .A2(\w[2][5] ),
    .A3(\w[6][5] ),
    .S0(net478),
    .S1(net486),
    .X(_07601_));
 sky130_fd_sc_hd__mux4_2 _19301_ (.A0(\w[8][5] ),
    .A1(\w[12][5] ),
    .A2(\w[10][5] ),
    .A3(\w[14][5] ),
    .S0(net478),
    .S1(net486),
    .X(_07602_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1020 ();
 sky130_fd_sc_hd__mux4_2 _19303_ (.A0(\w[16][5] ),
    .A1(\w[20][5] ),
    .A2(\w[18][5] ),
    .A3(\w[22][5] ),
    .S0(net478),
    .S1(net486),
    .X(_07604_));
 sky130_fd_sc_hd__mux4_2 _19304_ (.A0(\w[24][5] ),
    .A1(\w[28][5] ),
    .A2(\w[26][5] ),
    .A3(\w[30][5] ),
    .S0(net478),
    .S1(net486),
    .X(_07605_));
 sky130_fd_sc_hd__mux4_2 _19305_ (.A0(_07601_),
    .A1(_07602_),
    .A2(_07604_),
    .A3(_07605_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07606_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1019 ();
 sky130_fd_sc_hd__mux4_2 _19307_ (.A0(\w[32][5] ),
    .A1(\w[36][5] ),
    .A2(\w[34][5] ),
    .A3(\w[38][5] ),
    .S0(net478),
    .S1(net486),
    .X(_07608_));
 sky130_fd_sc_hd__mux4_2 _19308_ (.A0(\w[40][5] ),
    .A1(\w[44][5] ),
    .A2(\w[42][5] ),
    .A3(\w[46][5] ),
    .S0(net478),
    .S1(net486),
    .X(_07609_));
 sky130_fd_sc_hd__mux4_2 _19309_ (.A0(\w[48][5] ),
    .A1(\w[52][5] ),
    .A2(\w[50][5] ),
    .A3(\w[54][5] ),
    .S0(net478),
    .S1(net486),
    .X(_07610_));
 sky130_fd_sc_hd__mux4_2 _19310_ (.A0(\w[56][5] ),
    .A1(\w[60][5] ),
    .A2(\w[58][5] ),
    .A3(\w[62][5] ),
    .S0(net485),
    .S1(net486),
    .X(_07611_));
 sky130_fd_sc_hd__mux4_2 _19311_ (.A0(_07608_),
    .A1(_07609_),
    .A2(_07610_),
    .A3(_07611_),
    .S0(net546),
    .S1(net474),
    .X(_07612_));
 sky130_fd_sc_hd__mux2i_4 _19312_ (.A0(_07606_),
    .A1(_07612_),
    .S(net545),
    .Y(_11621_));
 sky130_fd_sc_hd__mux4_2 _19313_ (.A0(\w[0][6] ),
    .A1(\w[4][6] ),
    .A2(\w[2][6] ),
    .A3(\w[6][6] ),
    .S0(net485),
    .S1(net486),
    .X(_07613_));
 sky130_fd_sc_hd__mux4_2 _19314_ (.A0(\w[8][6] ),
    .A1(\w[12][6] ),
    .A2(\w[10][6] ),
    .A3(\w[14][6] ),
    .S0(net485),
    .S1(net486),
    .X(_07614_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1018 ();
 sky130_fd_sc_hd__mux4_2 _19316_ (.A0(\w[16][6] ),
    .A1(\w[20][6] ),
    .A2(\w[18][6] ),
    .A3(\w[22][6] ),
    .S0(net485),
    .S1(net486),
    .X(_07616_));
 sky130_fd_sc_hd__mux4_2 _19317_ (.A0(\w[24][6] ),
    .A1(\w[28][6] ),
    .A2(\w[26][6] ),
    .A3(\w[30][6] ),
    .S0(net485),
    .S1(net486),
    .X(_07617_));
 sky130_fd_sc_hd__mux4_2 _19318_ (.A0(_07613_),
    .A1(_07614_),
    .A2(_07616_),
    .A3(_07617_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07618_));
 sky130_fd_sc_hd__mux4_2 _19319_ (.A0(\w[32][6] ),
    .A1(\w[36][6] ),
    .A2(\w[34][6] ),
    .A3(\w[38][6] ),
    .S0(\count16_1[2] ),
    .S1(net491),
    .X(_07619_));
 sky130_fd_sc_hd__mux4_2 _19320_ (.A0(\w[40][6] ),
    .A1(\w[44][6] ),
    .A2(\w[42][6] ),
    .A3(\w[46][6] ),
    .S0(\count16_1[2] ),
    .S1(net491),
    .X(_07620_));
 sky130_fd_sc_hd__mux4_2 _19321_ (.A0(\w[48][6] ),
    .A1(\w[52][6] ),
    .A2(\w[50][6] ),
    .A3(\w[54][6] ),
    .S0(\count16_1[2] ),
    .S1(net491),
    .X(_07621_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1017 ();
 sky130_fd_sc_hd__mux4_2 _19323_ (.A0(\w[56][6] ),
    .A1(\w[60][6] ),
    .A2(\w[58][6] ),
    .A3(\w[62][6] ),
    .S0(\count16_1[2] ),
    .S1(net491),
    .X(_07623_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1016 ();
 sky130_fd_sc_hd__mux4_2 _19325_ (.A0(_07619_),
    .A1(_07620_),
    .A2(_07621_),
    .A3(_07623_),
    .S0(net546),
    .S1(net474),
    .X(_07625_));
 sky130_fd_sc_hd__mux2i_4 _19326_ (.A0(_07618_),
    .A1(_07625_),
    .S(net545),
    .Y(_11629_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1015 ();
 sky130_fd_sc_hd__mux4_2 _19328_ (.A0(\w[0][7] ),
    .A1(\w[4][7] ),
    .A2(\w[2][7] ),
    .A3(\w[6][7] ),
    .S0(net478),
    .S1(net486),
    .X(_07627_));
 sky130_fd_sc_hd__mux4_2 _19329_ (.A0(\w[8][7] ),
    .A1(\w[12][7] ),
    .A2(\w[10][7] ),
    .A3(\w[14][7] ),
    .S0(net478),
    .S1(net486),
    .X(_07628_));
 sky130_fd_sc_hd__mux4_2 _19330_ (.A0(\w[16][7] ),
    .A1(\w[20][7] ),
    .A2(\w[18][7] ),
    .A3(\w[22][7] ),
    .S0(net478),
    .S1(net486),
    .X(_07629_));
 sky130_fd_sc_hd__mux4_2 _19331_ (.A0(\w[24][7] ),
    .A1(\w[28][7] ),
    .A2(\w[26][7] ),
    .A3(\w[30][7] ),
    .S0(net478),
    .S1(net486),
    .X(_07630_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1014 ();
 sky130_fd_sc_hd__mux4_2 _19333_ (.A0(_07627_),
    .A1(_07628_),
    .A2(_07629_),
    .A3(_07630_),
    .S0(net546),
    .S1(net474),
    .X(_07632_));
 sky130_fd_sc_hd__mux4_2 _19334_ (.A0(\w[32][7] ),
    .A1(\w[36][7] ),
    .A2(\w[34][7] ),
    .A3(\w[38][7] ),
    .S0(\count16_1[2] ),
    .S1(net491),
    .X(_07633_));
 sky130_fd_sc_hd__mux4_2 _19335_ (.A0(\w[40][7] ),
    .A1(\w[44][7] ),
    .A2(\w[42][7] ),
    .A3(\w[46][7] ),
    .S0(\count16_1[2] ),
    .S1(net491),
    .X(_07634_));
 sky130_fd_sc_hd__mux4_2 _19336_ (.A0(\w[48][7] ),
    .A1(\w[52][7] ),
    .A2(\w[50][7] ),
    .A3(\w[54][7] ),
    .S0(\count16_1[2] ),
    .S1(net491),
    .X(_07635_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1013 ();
 sky130_fd_sc_hd__mux4_2 _19338_ (.A0(\w[56][7] ),
    .A1(\w[60][7] ),
    .A2(\w[58][7] ),
    .A3(\w[62][7] ),
    .S0(\count16_1[2] ),
    .S1(net491),
    .X(_07637_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1012 ();
 sky130_fd_sc_hd__mux4_2 _19340_ (.A0(_07633_),
    .A1(_07634_),
    .A2(_07635_),
    .A3(_07637_),
    .S0(net546),
    .S1(net474),
    .X(_07639_));
 sky130_fd_sc_hd__mux2i_4 _19341_ (.A0(_07632_),
    .A1(_07639_),
    .S(net545),
    .Y(_11637_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1011 ();
 sky130_fd_sc_hd__mux4_2 _19343_ (.A0(\w[0][8] ),
    .A1(\w[4][8] ),
    .A2(\w[2][8] ),
    .A3(\w[6][8] ),
    .S0(net480),
    .S1(net487),
    .X(_07641_));
 sky130_fd_sc_hd__mux4_2 _19344_ (.A0(\w[8][8] ),
    .A1(\w[12][8] ),
    .A2(\w[10][8] ),
    .A3(\w[14][8] ),
    .S0(net480),
    .S1(net487),
    .X(_07642_));
 sky130_fd_sc_hd__mux4_2 _19345_ (.A0(\w[16][8] ),
    .A1(\w[20][8] ),
    .A2(\w[18][8] ),
    .A3(\w[22][8] ),
    .S0(net480),
    .S1(net487),
    .X(_07643_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1010 ();
 sky130_fd_sc_hd__mux4_2 _19347_ (.A0(\w[24][8] ),
    .A1(\w[28][8] ),
    .A2(\w[26][8] ),
    .A3(\w[30][8] ),
    .S0(net480),
    .S1(net487),
    .X(_07645_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1009 ();
 sky130_fd_sc_hd__mux4_2 _19349_ (.A0(_07641_),
    .A1(_07642_),
    .A2(_07643_),
    .A3(_07645_),
    .S0(net476),
    .S1(net475),
    .X(_07647_));
 sky130_fd_sc_hd__mux4_2 _19350_ (.A0(\w[32][8] ),
    .A1(\w[36][8] ),
    .A2(\w[34][8] ),
    .A3(\w[38][8] ),
    .S0(net480),
    .S1(net489),
    .X(_07648_));
 sky130_fd_sc_hd__mux4_2 _19351_ (.A0(\w[40][8] ),
    .A1(\w[44][8] ),
    .A2(\w[42][8] ),
    .A3(\w[46][8] ),
    .S0(net480),
    .S1(net489),
    .X(_07649_));
 sky130_fd_sc_hd__mux4_2 _19352_ (.A0(\w[48][8] ),
    .A1(\w[52][8] ),
    .A2(\w[50][8] ),
    .A3(\w[54][8] ),
    .S0(net480),
    .S1(net489),
    .X(_07650_));
 sky130_fd_sc_hd__mux4_2 _19353_ (.A0(\w[56][8] ),
    .A1(\w[60][8] ),
    .A2(\w[58][8] ),
    .A3(\w[62][8] ),
    .S0(net480),
    .S1(net489),
    .X(_07651_));
 sky130_fd_sc_hd__mux4_2 _19354_ (.A0(_07648_),
    .A1(_07649_),
    .A2(_07650_),
    .A3(_07651_),
    .S0(net477),
    .S1(net475),
    .X(_07652_));
 sky130_fd_sc_hd__mux2i_4 _19355_ (.A0(_07647_),
    .A1(_07652_),
    .S(net472),
    .Y(_11645_));
 sky130_fd_sc_hd__mux4_2 _19356_ (.A0(\w[0][9] ),
    .A1(\w[4][9] ),
    .A2(\w[2][9] ),
    .A3(\w[6][9] ),
    .S0(net479),
    .S1(net489),
    .X(_07653_));
 sky130_fd_sc_hd__mux4_2 _19357_ (.A0(\w[8][9] ),
    .A1(\w[12][9] ),
    .A2(\w[10][9] ),
    .A3(\w[14][9] ),
    .S0(net479),
    .S1(net489),
    .X(_07654_));
 sky130_fd_sc_hd__mux4_2 _19358_ (.A0(\w[16][9] ),
    .A1(\w[20][9] ),
    .A2(\w[18][9] ),
    .A3(\w[22][9] ),
    .S0(net479),
    .S1(net489),
    .X(_07655_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1008 ();
 sky130_fd_sc_hd__mux4_2 _19360_ (.A0(\w[24][9] ),
    .A1(\w[28][9] ),
    .A2(\w[26][9] ),
    .A3(\w[30][9] ),
    .S0(net479),
    .S1(net489),
    .X(_07657_));
 sky130_fd_sc_hd__mux4_2 _19361_ (.A0(_07653_),
    .A1(_07654_),
    .A2(_07655_),
    .A3(_07657_),
    .S0(net477),
    .S1(net475),
    .X(_07658_));
 sky130_fd_sc_hd__mux4_2 _19362_ (.A0(\w[32][9] ),
    .A1(\w[36][9] ),
    .A2(\w[34][9] ),
    .A3(\w[38][9] ),
    .S0(net480),
    .S1(net489),
    .X(_07659_));
 sky130_fd_sc_hd__mux4_2 _19363_ (.A0(\w[40][9] ),
    .A1(\w[44][9] ),
    .A2(\w[42][9] ),
    .A3(\w[46][9] ),
    .S0(net480),
    .S1(net489),
    .X(_07660_));
 sky130_fd_sc_hd__mux4_2 _19364_ (.A0(\w[48][9] ),
    .A1(\w[52][9] ),
    .A2(\w[50][9] ),
    .A3(\w[54][9] ),
    .S0(net480),
    .S1(net489),
    .X(_07661_));
 sky130_fd_sc_hd__mux4_2 _19365_ (.A0(\w[56][9] ),
    .A1(\w[60][9] ),
    .A2(\w[58][9] ),
    .A3(\w[62][9] ),
    .S0(net480),
    .S1(net489),
    .X(_07662_));
 sky130_fd_sc_hd__mux4_2 _19366_ (.A0(_07659_),
    .A1(_07660_),
    .A2(_07661_),
    .A3(_07662_),
    .S0(net477),
    .S1(net475),
    .X(_07663_));
 sky130_fd_sc_hd__mux2i_4 _19367_ (.A0(_07658_),
    .A1(_07663_),
    .S(net472),
    .Y(_11653_));
 sky130_fd_sc_hd__mux4_2 _19368_ (.A0(\w[0][10] ),
    .A1(\w[4][10] ),
    .A2(\w[2][10] ),
    .A3(\w[6][10] ),
    .S0(net479),
    .S1(net489),
    .X(_07664_));
 sky130_fd_sc_hd__mux4_2 _19369_ (.A0(\w[8][10] ),
    .A1(\w[12][10] ),
    .A2(\w[10][10] ),
    .A3(\w[14][10] ),
    .S0(net479),
    .S1(net489),
    .X(_07665_));
 sky130_fd_sc_hd__mux4_2 _19370_ (.A0(\w[16][10] ),
    .A1(\w[20][10] ),
    .A2(\w[18][10] ),
    .A3(\w[22][10] ),
    .S0(net479),
    .S1(net489),
    .X(_07666_));
 sky130_fd_sc_hd__mux4_2 _19371_ (.A0(\w[24][10] ),
    .A1(\w[28][10] ),
    .A2(\w[26][10] ),
    .A3(\w[30][10] ),
    .S0(net479),
    .S1(net489),
    .X(_07667_));
 sky130_fd_sc_hd__mux4_2 _19372_ (.A0(_07664_),
    .A1(_07665_),
    .A2(_07666_),
    .A3(_07667_),
    .S0(net477),
    .S1(net475),
    .X(_07668_));
 sky130_fd_sc_hd__mux4_2 _19373_ (.A0(\w[32][10] ),
    .A1(\w[36][10] ),
    .A2(\w[34][10] ),
    .A3(\w[38][10] ),
    .S0(net484),
    .S1(net490),
    .X(_07669_));
 sky130_fd_sc_hd__mux4_2 _19374_ (.A0(\w[40][10] ),
    .A1(\w[44][10] ),
    .A2(\w[42][10] ),
    .A3(\w[46][10] ),
    .S0(net484),
    .S1(net490),
    .X(_07670_));
 sky130_fd_sc_hd__mux4_2 _19375_ (.A0(\w[48][10] ),
    .A1(\w[52][10] ),
    .A2(\w[50][10] ),
    .A3(\w[54][10] ),
    .S0(net484),
    .S1(net490),
    .X(_07671_));
 sky130_fd_sc_hd__mux4_2 _19376_ (.A0(\w[56][10] ),
    .A1(\w[60][10] ),
    .A2(\w[58][10] ),
    .A3(\w[62][10] ),
    .S0(net484),
    .S1(net490),
    .X(_07672_));
 sky130_fd_sc_hd__mux4_2 _19377_ (.A0(_07669_),
    .A1(_07670_),
    .A2(_07671_),
    .A3(_07672_),
    .S0(net477),
    .S1(net475),
    .X(_07673_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1007 ();
 sky130_fd_sc_hd__mux2i_4 _19379_ (.A0(_07668_),
    .A1(_07673_),
    .S(net472),
    .Y(_11661_));
 sky130_fd_sc_hd__mux4_2 _19380_ (.A0(\w[0][11] ),
    .A1(\w[4][11] ),
    .A2(\w[2][11] ),
    .A3(\w[6][11] ),
    .S0(net480),
    .S1(net487),
    .X(_07675_));
 sky130_fd_sc_hd__mux4_2 _19381_ (.A0(\w[8][11] ),
    .A1(\w[12][11] ),
    .A2(\w[10][11] ),
    .A3(\w[14][11] ),
    .S0(net482),
    .S1(net487),
    .X(_07676_));
 sky130_fd_sc_hd__mux4_2 _19382_ (.A0(\w[16][11] ),
    .A1(\w[20][11] ),
    .A2(\w[18][11] ),
    .A3(\w[22][11] ),
    .S0(net480),
    .S1(net487),
    .X(_07677_));
 sky130_fd_sc_hd__mux4_2 _19383_ (.A0(\w[24][11] ),
    .A1(\w[28][11] ),
    .A2(\w[26][11] ),
    .A3(\w[30][11] ),
    .S0(net480),
    .S1(net487),
    .X(_07678_));
 sky130_fd_sc_hd__mux4_2 _19384_ (.A0(_07675_),
    .A1(_07676_),
    .A2(_07677_),
    .A3(_07678_),
    .S0(net476),
    .S1(net475),
    .X(_07679_));
 sky130_fd_sc_hd__mux4_2 _19385_ (.A0(\w[32][11] ),
    .A1(\w[36][11] ),
    .A2(\w[34][11] ),
    .A3(\w[38][11] ),
    .S0(net484),
    .S1(net490),
    .X(_07680_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1006 ();
 sky130_fd_sc_hd__mux4_2 _19387_ (.A0(\w[40][11] ),
    .A1(\w[44][11] ),
    .A2(\w[42][11] ),
    .A3(\w[46][11] ),
    .S0(net484),
    .S1(net490),
    .X(_07682_));
 sky130_fd_sc_hd__mux4_2 _19388_ (.A0(\w[48][11] ),
    .A1(\w[52][11] ),
    .A2(\w[50][11] ),
    .A3(\w[54][11] ),
    .S0(net484),
    .S1(net490),
    .X(_07683_));
 sky130_fd_sc_hd__mux4_2 _19389_ (.A0(\w[56][11] ),
    .A1(\w[60][11] ),
    .A2(\w[58][11] ),
    .A3(\w[62][11] ),
    .S0(net484),
    .S1(net490),
    .X(_07684_));
 sky130_fd_sc_hd__mux4_2 _19390_ (.A0(_07680_),
    .A1(_07682_),
    .A2(_07683_),
    .A3(_07684_),
    .S0(net477),
    .S1(\count16_1[4] ),
    .X(_07685_));
 sky130_fd_sc_hd__mux2i_2 _19391_ (.A0(_07679_),
    .A1(_07685_),
    .S(net472),
    .Y(_11669_));
 sky130_fd_sc_hd__mux4_2 _19392_ (.A0(\w[0][12] ),
    .A1(\w[4][12] ),
    .A2(\w[2][12] ),
    .A3(\w[6][12] ),
    .S0(net483),
    .S1(net491),
    .X(_07686_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1005 ();
 sky130_fd_sc_hd__mux4_2 _19394_ (.A0(\w[8][12] ),
    .A1(\w[12][12] ),
    .A2(\w[10][12] ),
    .A3(\w[14][12] ),
    .S0(net483),
    .S1(net491),
    .X(_07688_));
 sky130_fd_sc_hd__mux4_2 _19395_ (.A0(\w[16][12] ),
    .A1(\w[20][12] ),
    .A2(\w[18][12] ),
    .A3(\w[22][12] ),
    .S0(net483),
    .S1(net491),
    .X(_07689_));
 sky130_fd_sc_hd__mux4_2 _19396_ (.A0(\w[24][12] ),
    .A1(\w[28][12] ),
    .A2(\w[26][12] ),
    .A3(\w[30][12] ),
    .S0(net483),
    .S1(net491),
    .X(_07690_));
 sky130_fd_sc_hd__mux4_2 _19397_ (.A0(_07686_),
    .A1(_07688_),
    .A2(_07689_),
    .A3(_07690_),
    .S0(net476),
    .S1(net474),
    .X(_07691_));
 sky130_fd_sc_hd__mux4_2 _19398_ (.A0(\w[32][12] ),
    .A1(\w[36][12] ),
    .A2(\w[34][12] ),
    .A3(\w[38][12] ),
    .S0(net483),
    .S1(net491),
    .X(_07692_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1004 ();
 sky130_fd_sc_hd__mux4_2 _19400_ (.A0(\w[40][12] ),
    .A1(\w[44][12] ),
    .A2(\w[42][12] ),
    .A3(\w[46][12] ),
    .S0(net483),
    .S1(net488),
    .X(_07694_));
 sky130_fd_sc_hd__mux4_2 _19401_ (.A0(\w[48][12] ),
    .A1(\w[52][12] ),
    .A2(\w[50][12] ),
    .A3(\w[54][12] ),
    .S0(net483),
    .S1(net491),
    .X(_07695_));
 sky130_fd_sc_hd__mux4_2 _19402_ (.A0(\w[56][12] ),
    .A1(\w[60][12] ),
    .A2(\w[58][12] ),
    .A3(\w[62][12] ),
    .S0(net483),
    .S1(net491),
    .X(_07696_));
 sky130_fd_sc_hd__mux4_2 _19403_ (.A0(_07692_),
    .A1(_07694_),
    .A2(_07695_),
    .A3(_07696_),
    .S0(net476),
    .S1(net474),
    .X(_07697_));
 sky130_fd_sc_hd__mux2i_4 _19404_ (.A0(_07691_),
    .A1(_07697_),
    .S(net545),
    .Y(_11677_));
 sky130_fd_sc_hd__mux4_2 _19405_ (.A0(\w[0][13] ),
    .A1(\w[4][13] ),
    .A2(\w[2][13] ),
    .A3(\w[6][13] ),
    .S0(net482),
    .S1(net487),
    .X(_07698_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1003 ();
 sky130_fd_sc_hd__mux4_2 _19407_ (.A0(\w[8][13] ),
    .A1(\w[12][13] ),
    .A2(\w[10][13] ),
    .A3(\w[14][13] ),
    .S0(net482),
    .S1(net487),
    .X(_07700_));
 sky130_fd_sc_hd__mux4_2 _19408_ (.A0(\w[16][13] ),
    .A1(\w[20][13] ),
    .A2(\w[18][13] ),
    .A3(\w[22][13] ),
    .S0(net482),
    .S1(net487),
    .X(_07701_));
 sky130_fd_sc_hd__mux4_2 _19409_ (.A0(\w[24][13] ),
    .A1(\w[28][13] ),
    .A2(\w[26][13] ),
    .A3(\w[30][13] ),
    .S0(net482),
    .S1(net487),
    .X(_07702_));
 sky130_fd_sc_hd__mux4_2 _19410_ (.A0(_07698_),
    .A1(_07700_),
    .A2(_07701_),
    .A3(_07702_),
    .S0(net476),
    .S1(net474),
    .X(_07703_));
 sky130_fd_sc_hd__mux4_2 _19411_ (.A0(\w[32][13] ),
    .A1(\w[36][13] ),
    .A2(\w[34][13] ),
    .A3(\w[38][13] ),
    .S0(net482),
    .S1(net489),
    .X(_07704_));
 sky130_fd_sc_hd__mux4_2 _19412_ (.A0(\w[40][13] ),
    .A1(\w[44][13] ),
    .A2(\w[42][13] ),
    .A3(\w[46][13] ),
    .S0(net482),
    .S1(net490),
    .X(_07705_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1002 ();
 sky130_fd_sc_hd__mux4_2 _19414_ (.A0(\w[48][13] ),
    .A1(\w[52][13] ),
    .A2(\w[50][13] ),
    .A3(\w[54][13] ),
    .S0(net483),
    .S1(net490),
    .X(_07707_));
 sky130_fd_sc_hd__mux4_2 _19415_ (.A0(\w[56][13] ),
    .A1(\w[60][13] ),
    .A2(\w[58][13] ),
    .A3(\w[62][13] ),
    .S0(\count16_1[2] ),
    .S1(net490),
    .X(_07708_));
 sky130_fd_sc_hd__mux4_2 _19416_ (.A0(_07704_),
    .A1(_07705_),
    .A2(_07707_),
    .A3(_07708_),
    .S0(net546),
    .S1(net474),
    .X(_07709_));
 sky130_fd_sc_hd__mux2i_2 _19417_ (.A0(_07703_),
    .A1(_07709_),
    .S(net473),
    .Y(_11685_));
 sky130_fd_sc_hd__mux4_2 _19418_ (.A0(\w[0][14] ),
    .A1(\w[4][14] ),
    .A2(\w[2][14] ),
    .A3(\w[6][14] ),
    .S0(net483),
    .S1(net491),
    .X(_07710_));
 sky130_fd_sc_hd__mux4_2 _19419_ (.A0(\w[8][14] ),
    .A1(\w[12][14] ),
    .A2(\w[10][14] ),
    .A3(\w[14][14] ),
    .S0(net483),
    .S1(net491),
    .X(_07711_));
 sky130_fd_sc_hd__mux4_2 _19420_ (.A0(\w[16][14] ),
    .A1(\w[20][14] ),
    .A2(\w[18][14] ),
    .A3(\w[22][14] ),
    .S0(net483),
    .S1(net491),
    .X(_07712_));
 sky130_fd_sc_hd__mux4_2 _19421_ (.A0(\w[24][14] ),
    .A1(\w[28][14] ),
    .A2(\w[26][14] ),
    .A3(\w[30][14] ),
    .S0(net483),
    .S1(net491),
    .X(_07713_));
 sky130_fd_sc_hd__mux4_2 _19422_ (.A0(_07710_),
    .A1(_07711_),
    .A2(_07712_),
    .A3(_07713_),
    .S0(net476),
    .S1(net474),
    .X(_07714_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1001 ();
 sky130_fd_sc_hd__mux4_2 _19424_ (.A0(\w[32][14] ),
    .A1(\w[36][14] ),
    .A2(\w[34][14] ),
    .A3(\w[38][14] ),
    .S0(net481),
    .S1(net489),
    .X(_07716_));
 sky130_fd_sc_hd__mux4_2 _19425_ (.A0(\w[40][14] ),
    .A1(\w[44][14] ),
    .A2(\w[42][14] ),
    .A3(\w[46][14] ),
    .S0(net481),
    .S1(net489),
    .X(_07717_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1000 ();
 sky130_fd_sc_hd__mux4_2 _19427_ (.A0(\w[48][14] ),
    .A1(\w[52][14] ),
    .A2(\w[50][14] ),
    .A3(\w[54][14] ),
    .S0(net481),
    .S1(net489),
    .X(_07719_));
 sky130_fd_sc_hd__mux4_2 _19428_ (.A0(\w[56][14] ),
    .A1(\w[60][14] ),
    .A2(\w[58][14] ),
    .A3(\w[62][14] ),
    .S0(net481),
    .S1(net489),
    .X(_07720_));
 sky130_fd_sc_hd__mux4_2 _19429_ (.A0(_07716_),
    .A1(_07717_),
    .A2(_07719_),
    .A3(_07720_),
    .S0(net476),
    .S1(net474),
    .X(_07721_));
 sky130_fd_sc_hd__mux2i_4 _19430_ (.A0(_07714_),
    .A1(_07721_),
    .S(net473),
    .Y(_11693_));
 sky130_fd_sc_hd__mux4_2 _19431_ (.A0(\w[0][15] ),
    .A1(\w[4][15] ),
    .A2(\w[2][15] ),
    .A3(\w[6][15] ),
    .S0(net485),
    .S1(net486),
    .X(_07722_));
 sky130_fd_sc_hd__mux4_2 _19432_ (.A0(\w[8][15] ),
    .A1(\w[12][15] ),
    .A2(\w[10][15] ),
    .A3(\w[14][15] ),
    .S0(net485),
    .S1(net486),
    .X(_07723_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_999 ();
 sky130_fd_sc_hd__mux4_2 _19434_ (.A0(\w[16][15] ),
    .A1(\w[20][15] ),
    .A2(\w[18][15] ),
    .A3(\w[22][15] ),
    .S0(net485),
    .S1(net486),
    .X(_07725_));
 sky130_fd_sc_hd__mux4_2 _19435_ (.A0(\w[24][15] ),
    .A1(\w[28][15] ),
    .A2(\w[26][15] ),
    .A3(\w[30][15] ),
    .S0(net485),
    .S1(net486),
    .X(_07726_));
 sky130_fd_sc_hd__mux4_2 _19436_ (.A0(_07722_),
    .A1(_07723_),
    .A2(_07725_),
    .A3(_07726_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07727_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_998 ();
 sky130_fd_sc_hd__mux4_2 _19438_ (.A0(\w[32][15] ),
    .A1(\w[36][15] ),
    .A2(\w[34][15] ),
    .A3(\w[38][15] ),
    .S0(net485),
    .S1(net486),
    .X(_07729_));
 sky130_fd_sc_hd__mux4_2 _19439_ (.A0(\w[40][15] ),
    .A1(\w[44][15] ),
    .A2(\w[42][15] ),
    .A3(\w[46][15] ),
    .S0(net485),
    .S1(net486),
    .X(_07730_));
 sky130_fd_sc_hd__mux4_2 _19440_ (.A0(\w[48][15] ),
    .A1(\w[52][15] ),
    .A2(\w[50][15] ),
    .A3(\w[54][15] ),
    .S0(net485),
    .S1(net486),
    .X(_07731_));
 sky130_fd_sc_hd__mux4_2 _19441_ (.A0(\w[56][15] ),
    .A1(\w[60][15] ),
    .A2(\w[58][15] ),
    .A3(\w[62][15] ),
    .S0(net485),
    .S1(net486),
    .X(_07732_));
 sky130_fd_sc_hd__mux4_2 _19442_ (.A0(_07729_),
    .A1(_07730_),
    .A2(_07731_),
    .A3(_07732_),
    .S0(net546),
    .S1(net474),
    .X(_07733_));
 sky130_fd_sc_hd__mux2i_4 _19443_ (.A0(_07727_),
    .A1(_07733_),
    .S(net545),
    .Y(_11701_));
 sky130_fd_sc_hd__mux4_2 _19444_ (.A0(\w[0][16] ),
    .A1(\w[4][16] ),
    .A2(\w[2][16] ),
    .A3(\w[6][16] ),
    .S0(net485),
    .S1(net486),
    .X(_07734_));
 sky130_fd_sc_hd__mux4_2 _19445_ (.A0(\w[8][16] ),
    .A1(\w[12][16] ),
    .A2(\w[10][16] ),
    .A3(\w[14][16] ),
    .S0(net485),
    .S1(\count16_1[1] ),
    .X(_07735_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_997 ();
 sky130_fd_sc_hd__mux4_2 _19447_ (.A0(\w[16][16] ),
    .A1(\w[20][16] ),
    .A2(\w[18][16] ),
    .A3(\w[22][16] ),
    .S0(net485),
    .S1(\count16_1[1] ),
    .X(_07737_));
 sky130_fd_sc_hd__mux4_2 _19448_ (.A0(\w[24][16] ),
    .A1(\w[28][16] ),
    .A2(\w[26][16] ),
    .A3(\w[30][16] ),
    .S0(net485),
    .S1(\count16_1[1] ),
    .X(_07738_));
 sky130_fd_sc_hd__mux4_2 _19449_ (.A0(_07734_),
    .A1(_07735_),
    .A2(_07737_),
    .A3(_07738_),
    .S0(\count16_1[3] ),
    .S1(\count16_1[4] ),
    .X(_07739_));
 sky130_fd_sc_hd__mux4_2 _19450_ (.A0(\w[32][16] ),
    .A1(\w[36][16] ),
    .A2(\w[34][16] ),
    .A3(\w[38][16] ),
    .S0(\count16_1[2] ),
    .S1(net490),
    .X(_07740_));
 sky130_fd_sc_hd__mux4_2 _19451_ (.A0(\w[40][16] ),
    .A1(\w[44][16] ),
    .A2(\w[42][16] ),
    .A3(\w[46][16] ),
    .S0(\count16_1[2] ),
    .S1(net490),
    .X(_07741_));
 sky130_fd_sc_hd__mux4_2 _19452_ (.A0(\w[48][16] ),
    .A1(\w[52][16] ),
    .A2(\w[50][16] ),
    .A3(\w[54][16] ),
    .S0(\count16_1[2] ),
    .S1(net490),
    .X(_07742_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_996 ();
 sky130_fd_sc_hd__mux4_2 _19454_ (.A0(\w[56][16] ),
    .A1(\w[60][16] ),
    .A2(\w[58][16] ),
    .A3(\w[62][16] ),
    .S0(\count16_1[2] ),
    .S1(net490),
    .X(_07744_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_995 ();
 sky130_fd_sc_hd__mux4_2 _19456_ (.A0(_07740_),
    .A1(_07741_),
    .A2(_07742_),
    .A3(_07744_),
    .S0(net477),
    .S1(\count16_1[4] ),
    .X(_07746_));
 sky130_fd_sc_hd__mux2i_2 _19457_ (.A0(_07739_),
    .A1(_07746_),
    .S(net545),
    .Y(_11709_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_994 ();
 sky130_fd_sc_hd__mux4_2 _19459_ (.A0(\w[0][17] ),
    .A1(\w[4][17] ),
    .A2(\w[2][17] ),
    .A3(\w[6][17] ),
    .S0(net482),
    .S1(net487),
    .X(_07748_));
 sky130_fd_sc_hd__mux4_2 _19460_ (.A0(\w[8][17] ),
    .A1(\w[12][17] ),
    .A2(\w[10][17] ),
    .A3(\w[14][17] ),
    .S0(net482),
    .S1(net487),
    .X(_07749_));
 sky130_fd_sc_hd__mux4_2 _19461_ (.A0(\w[16][17] ),
    .A1(\w[20][17] ),
    .A2(\w[18][17] ),
    .A3(\w[22][17] ),
    .S0(net482),
    .S1(net487),
    .X(_07750_));
 sky130_fd_sc_hd__mux4_2 _19462_ (.A0(\w[24][17] ),
    .A1(\w[28][17] ),
    .A2(\w[26][17] ),
    .A3(\w[30][17] ),
    .S0(net482),
    .S1(net487),
    .X(_07751_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_993 ();
 sky130_fd_sc_hd__mux4_2 _19464_ (.A0(_07748_),
    .A1(_07749_),
    .A2(_07750_),
    .A3(_07751_),
    .S0(net476),
    .S1(net474),
    .X(_07753_));
 sky130_fd_sc_hd__mux4_2 _19465_ (.A0(\w[32][17] ),
    .A1(\w[36][17] ),
    .A2(\w[34][17] ),
    .A3(\w[38][17] ),
    .S0(net482),
    .S1(net488),
    .X(_07754_));
 sky130_fd_sc_hd__mux4_2 _19466_ (.A0(\w[40][17] ),
    .A1(\w[44][17] ),
    .A2(\w[42][17] ),
    .A3(\w[46][17] ),
    .S0(net482),
    .S1(net488),
    .X(_07755_));
 sky130_fd_sc_hd__mux4_2 _19467_ (.A0(\w[48][17] ),
    .A1(\w[52][17] ),
    .A2(\w[50][17] ),
    .A3(\w[54][17] ),
    .S0(net482),
    .S1(net488),
    .X(_07756_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_992 ();
 sky130_fd_sc_hd__mux4_2 _19469_ (.A0(\w[56][17] ),
    .A1(\w[60][17] ),
    .A2(\w[58][17] ),
    .A3(\w[62][17] ),
    .S0(net482),
    .S1(net488),
    .X(_07758_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_991 ();
 sky130_fd_sc_hd__mux4_2 _19471_ (.A0(_07754_),
    .A1(_07755_),
    .A2(_07756_),
    .A3(_07758_),
    .S0(net476),
    .S1(net474),
    .X(_07760_));
 sky130_fd_sc_hd__mux2i_4 _19472_ (.A0(_07753_),
    .A1(_07760_),
    .S(net473),
    .Y(_11717_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_990 ();
 sky130_fd_sc_hd__mux4_2 _19474_ (.A0(\w[0][18] ),
    .A1(\w[4][18] ),
    .A2(\w[2][18] ),
    .A3(\w[6][18] ),
    .S0(net484),
    .S1(net490),
    .X(_07762_));
 sky130_fd_sc_hd__mux4_2 _19475_ (.A0(\w[8][18] ),
    .A1(\w[12][18] ),
    .A2(\w[10][18] ),
    .A3(\w[14][18] ),
    .S0(net484),
    .S1(net490),
    .X(_07763_));
 sky130_fd_sc_hd__mux4_2 _19476_ (.A0(\w[16][18] ),
    .A1(\w[20][18] ),
    .A2(\w[18][18] ),
    .A3(\w[22][18] ),
    .S0(net484),
    .S1(net490),
    .X(_07764_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_989 ();
 sky130_fd_sc_hd__mux4_2 _19478_ (.A0(\w[24][18] ),
    .A1(\w[28][18] ),
    .A2(\w[26][18] ),
    .A3(\w[30][18] ),
    .S0(net484),
    .S1(net490),
    .X(_07766_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_988 ();
 sky130_fd_sc_hd__mux4_2 _19480_ (.A0(_07762_),
    .A1(_07763_),
    .A2(_07764_),
    .A3(_07766_),
    .S0(net477),
    .S1(net475),
    .X(_07768_));
 sky130_fd_sc_hd__mux4_2 _19481_ (.A0(\w[32][18] ),
    .A1(\w[36][18] ),
    .A2(\w[34][18] ),
    .A3(\w[38][18] ),
    .S0(net484),
    .S1(net490),
    .X(_07769_));
 sky130_fd_sc_hd__mux4_2 _19482_ (.A0(\w[40][18] ),
    .A1(\w[44][18] ),
    .A2(\w[42][18] ),
    .A3(\w[46][18] ),
    .S0(net484),
    .S1(net490),
    .X(_07770_));
 sky130_fd_sc_hd__mux4_2 _19483_ (.A0(\w[48][18] ),
    .A1(\w[52][18] ),
    .A2(\w[50][18] ),
    .A3(\w[54][18] ),
    .S0(net484),
    .S1(net490),
    .X(_07771_));
 sky130_fd_sc_hd__mux4_2 _19484_ (.A0(\w[56][18] ),
    .A1(\w[60][18] ),
    .A2(\w[58][18] ),
    .A3(\w[62][18] ),
    .S0(net484),
    .S1(net490),
    .X(_07772_));
 sky130_fd_sc_hd__mux4_2 _19485_ (.A0(_07769_),
    .A1(_07770_),
    .A2(_07771_),
    .A3(_07772_),
    .S0(net477),
    .S1(net475),
    .X(_07773_));
 sky130_fd_sc_hd__mux2i_2 _19486_ (.A0(_07768_),
    .A1(_07773_),
    .S(net472),
    .Y(_11725_));
 sky130_fd_sc_hd__mux4_2 _19487_ (.A0(\w[0][19] ),
    .A1(\w[4][19] ),
    .A2(\w[2][19] ),
    .A3(\w[6][19] ),
    .S0(net480),
    .S1(net487),
    .X(_07774_));
 sky130_fd_sc_hd__mux4_2 _19488_ (.A0(\w[8][19] ),
    .A1(\w[12][19] ),
    .A2(\w[10][19] ),
    .A3(\w[14][19] ),
    .S0(net480),
    .S1(net487),
    .X(_07775_));
 sky130_fd_sc_hd__mux4_2 _19489_ (.A0(\w[16][19] ),
    .A1(\w[20][19] ),
    .A2(\w[18][19] ),
    .A3(\w[22][19] ),
    .S0(net480),
    .S1(net487),
    .X(_07776_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_987 ();
 sky130_fd_sc_hd__mux4_2 _19491_ (.A0(\w[24][19] ),
    .A1(\w[28][19] ),
    .A2(\w[26][19] ),
    .A3(\w[30][19] ),
    .S0(net480),
    .S1(net487),
    .X(_07778_));
 sky130_fd_sc_hd__mux4_2 _19492_ (.A0(_07774_),
    .A1(_07775_),
    .A2(_07776_),
    .A3(_07778_),
    .S0(net476),
    .S1(net475),
    .X(_07779_));
 sky130_fd_sc_hd__mux4_2 _19493_ (.A0(\w[32][19] ),
    .A1(\w[36][19] ),
    .A2(\w[34][19] ),
    .A3(\w[38][19] ),
    .S0(net484),
    .S1(net490),
    .X(_07780_));
 sky130_fd_sc_hd__mux4_2 _19494_ (.A0(\w[40][19] ),
    .A1(\w[44][19] ),
    .A2(\w[42][19] ),
    .A3(\w[46][19] ),
    .S0(net484),
    .S1(net490),
    .X(_07781_));
 sky130_fd_sc_hd__mux4_2 _19495_ (.A0(\w[48][19] ),
    .A1(\w[52][19] ),
    .A2(\w[50][19] ),
    .A3(\w[54][19] ),
    .S0(net484),
    .S1(net490),
    .X(_07782_));
 sky130_fd_sc_hd__mux4_2 _19496_ (.A0(\w[56][19] ),
    .A1(\w[60][19] ),
    .A2(\w[58][19] ),
    .A3(\w[62][19] ),
    .S0(net484),
    .S1(net490),
    .X(_07783_));
 sky130_fd_sc_hd__mux4_2 _19497_ (.A0(_07780_),
    .A1(_07781_),
    .A2(_07782_),
    .A3(_07783_),
    .S0(net477),
    .S1(net475),
    .X(_07784_));
 sky130_fd_sc_hd__mux2i_4 _19498_ (.A0(_07779_),
    .A1(_07784_),
    .S(net472),
    .Y(_11733_));
 sky130_fd_sc_hd__mux4_2 _19499_ (.A0(\w[0][20] ),
    .A1(\w[4][20] ),
    .A2(\w[2][20] ),
    .A3(\w[6][20] ),
    .S0(net484),
    .S1(net490),
    .X(_07785_));
 sky130_fd_sc_hd__mux4_2 _19500_ (.A0(\w[8][20] ),
    .A1(\w[12][20] ),
    .A2(\w[10][20] ),
    .A3(\w[14][20] ),
    .S0(net484),
    .S1(net490),
    .X(_07786_));
 sky130_fd_sc_hd__mux4_2 _19501_ (.A0(\w[16][20] ),
    .A1(\w[20][20] ),
    .A2(\w[18][20] ),
    .A3(\w[22][20] ),
    .S0(net484),
    .S1(net490),
    .X(_07787_));
 sky130_fd_sc_hd__mux4_2 _19502_ (.A0(\w[24][20] ),
    .A1(\w[28][20] ),
    .A2(\w[26][20] ),
    .A3(\w[30][20] ),
    .S0(net484),
    .S1(net490),
    .X(_07788_));
 sky130_fd_sc_hd__mux4_2 _19503_ (.A0(_07785_),
    .A1(_07786_),
    .A2(_07787_),
    .A3(_07788_),
    .S0(net477),
    .S1(net475),
    .X(_07789_));
 sky130_fd_sc_hd__mux4_2 _19504_ (.A0(\w[32][20] ),
    .A1(\w[36][20] ),
    .A2(\w[34][20] ),
    .A3(\w[38][20] ),
    .S0(net484),
    .S1(net490),
    .X(_07790_));
 sky130_fd_sc_hd__mux4_2 _19505_ (.A0(\w[40][20] ),
    .A1(\w[44][20] ),
    .A2(\w[42][20] ),
    .A3(\w[46][20] ),
    .S0(net484),
    .S1(net490),
    .X(_07791_));
 sky130_fd_sc_hd__mux4_2 _19506_ (.A0(\w[48][20] ),
    .A1(\w[52][20] ),
    .A2(\w[50][20] ),
    .A3(\w[54][20] ),
    .S0(net484),
    .S1(net490),
    .X(_07792_));
 sky130_fd_sc_hd__mux4_2 _19507_ (.A0(\w[56][20] ),
    .A1(\w[60][20] ),
    .A2(\w[58][20] ),
    .A3(\w[62][20] ),
    .S0(net484),
    .S1(net490),
    .X(_07793_));
 sky130_fd_sc_hd__mux4_2 _19508_ (.A0(_07790_),
    .A1(_07791_),
    .A2(_07792_),
    .A3(_07793_),
    .S0(net477),
    .S1(net475),
    .X(_07794_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_986 ();
 sky130_fd_sc_hd__mux2i_4 _19510_ (.A0(_07789_),
    .A1(_07794_),
    .S(net472),
    .Y(_11741_));
 sky130_fd_sc_hd__mux4_2 _19511_ (.A0(\w[0][21] ),
    .A1(\w[4][21] ),
    .A2(\w[2][21] ),
    .A3(\w[6][21] ),
    .S0(net480),
    .S1(net488),
    .X(_07796_));
 sky130_fd_sc_hd__mux4_2 _19512_ (.A0(\w[8][21] ),
    .A1(\w[12][21] ),
    .A2(\w[10][21] ),
    .A3(\w[14][21] ),
    .S0(net480),
    .S1(net488),
    .X(_07797_));
 sky130_fd_sc_hd__mux4_2 _19513_ (.A0(\w[16][21] ),
    .A1(\w[20][21] ),
    .A2(\w[18][21] ),
    .A3(\w[22][21] ),
    .S0(net480),
    .S1(net488),
    .X(_07798_));
 sky130_fd_sc_hd__mux4_2 _19514_ (.A0(\w[24][21] ),
    .A1(\w[28][21] ),
    .A2(\w[26][21] ),
    .A3(\w[30][21] ),
    .S0(net480),
    .S1(net488),
    .X(_07799_));
 sky130_fd_sc_hd__mux4_2 _19515_ (.A0(_07796_),
    .A1(_07797_),
    .A2(_07798_),
    .A3(_07799_),
    .S0(net476),
    .S1(net475),
    .X(_07800_));
 sky130_fd_sc_hd__mux4_2 _19516_ (.A0(\w[32][21] ),
    .A1(\w[36][21] ),
    .A2(\w[34][21] ),
    .A3(\w[38][21] ),
    .S0(net481),
    .S1(net489),
    .X(_07801_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_985 ();
 sky130_fd_sc_hd__mux4_2 _19518_ (.A0(\w[40][21] ),
    .A1(\w[44][21] ),
    .A2(\w[42][21] ),
    .A3(\w[46][21] ),
    .S0(net481),
    .S1(net489),
    .X(_07803_));
 sky130_fd_sc_hd__mux4_2 _19519_ (.A0(\w[48][21] ),
    .A1(\w[52][21] ),
    .A2(\w[50][21] ),
    .A3(\w[54][21] ),
    .S0(net481),
    .S1(net489),
    .X(_07804_));
 sky130_fd_sc_hd__mux4_2 _19520_ (.A0(\w[56][21] ),
    .A1(\w[60][21] ),
    .A2(\w[58][21] ),
    .A3(\w[62][21] ),
    .S0(net481),
    .S1(net489),
    .X(_07805_));
 sky130_fd_sc_hd__mux4_2 _19521_ (.A0(_07801_),
    .A1(_07803_),
    .A2(_07804_),
    .A3(_07805_),
    .S0(net477),
    .S1(net475),
    .X(_07806_));
 sky130_fd_sc_hd__mux2i_2 _19522_ (.A0(_07800_),
    .A1(_07806_),
    .S(net472),
    .Y(_11749_));
 sky130_fd_sc_hd__mux4_2 _19523_ (.A0(\w[0][22] ),
    .A1(\w[4][22] ),
    .A2(\w[2][22] ),
    .A3(\w[6][22] ),
    .S0(net479),
    .S1(net489),
    .X(_07807_));
 sky130_fd_sc_hd__mux4_2 _19524_ (.A0(\w[8][22] ),
    .A1(\w[12][22] ),
    .A2(\w[10][22] ),
    .A3(\w[14][22] ),
    .S0(net480),
    .S1(net487),
    .X(_07808_));
 sky130_fd_sc_hd__mux4_2 _19525_ (.A0(\w[16][22] ),
    .A1(\w[20][22] ),
    .A2(\w[18][22] ),
    .A3(\w[22][22] ),
    .S0(net480),
    .S1(net487),
    .X(_07809_));
 sky130_fd_sc_hd__mux4_2 _19526_ (.A0(\w[24][22] ),
    .A1(\w[28][22] ),
    .A2(\w[26][22] ),
    .A3(\w[30][22] ),
    .S0(net480),
    .S1(net487),
    .X(_07810_));
 sky130_fd_sc_hd__mux4_2 _19527_ (.A0(_07807_),
    .A1(_07808_),
    .A2(_07809_),
    .A3(_07810_),
    .S0(net477),
    .S1(net475),
    .X(_07811_));
 sky130_fd_sc_hd__mux4_2 _19528_ (.A0(\w[32][22] ),
    .A1(\w[36][22] ),
    .A2(\w[34][22] ),
    .A3(\w[38][22] ),
    .S0(net479),
    .S1(net489),
    .X(_07812_));
 sky130_fd_sc_hd__mux4_2 _19529_ (.A0(\w[40][22] ),
    .A1(\w[44][22] ),
    .A2(\w[42][22] ),
    .A3(\w[46][22] ),
    .S0(net479),
    .S1(net489),
    .X(_07813_));
 sky130_fd_sc_hd__mux4_2 _19530_ (.A0(\w[48][22] ),
    .A1(\w[52][22] ),
    .A2(\w[50][22] ),
    .A3(\w[54][22] ),
    .S0(net479),
    .S1(net489),
    .X(_07814_));
 sky130_fd_sc_hd__mux4_2 _19531_ (.A0(\w[56][22] ),
    .A1(\w[60][22] ),
    .A2(\w[58][22] ),
    .A3(\w[62][22] ),
    .S0(net479),
    .S1(net489),
    .X(_07815_));
 sky130_fd_sc_hd__mux4_2 _19532_ (.A0(_07812_),
    .A1(_07813_),
    .A2(_07814_),
    .A3(_07815_),
    .S0(net477),
    .S1(net475),
    .X(_07816_));
 sky130_fd_sc_hd__mux2i_4 _19533_ (.A0(_07811_),
    .A1(_07816_),
    .S(net472),
    .Y(_11757_));
 sky130_fd_sc_hd__mux4_2 _19534_ (.A0(\w[0][23] ),
    .A1(\w[4][23] ),
    .A2(\w[2][23] ),
    .A3(\w[6][23] ),
    .S0(net483),
    .S1(net491),
    .X(_07817_));
 sky130_fd_sc_hd__mux4_2 _19535_ (.A0(\w[8][23] ),
    .A1(\w[12][23] ),
    .A2(\w[10][23] ),
    .A3(\w[14][23] ),
    .S0(net483),
    .S1(net491),
    .X(_07818_));
 sky130_fd_sc_hd__mux4_2 _19536_ (.A0(\w[16][23] ),
    .A1(\w[20][23] ),
    .A2(\w[18][23] ),
    .A3(\w[22][23] ),
    .S0(net483),
    .S1(net491),
    .X(_07819_));
 sky130_fd_sc_hd__mux4_2 _19537_ (.A0(\w[24][23] ),
    .A1(\w[28][23] ),
    .A2(\w[26][23] ),
    .A3(\w[30][23] ),
    .S0(net483),
    .S1(net491),
    .X(_07820_));
 sky130_fd_sc_hd__mux4_2 _19538_ (.A0(_07817_),
    .A1(_07818_),
    .A2(_07819_),
    .A3(_07820_),
    .S0(net476),
    .S1(net474),
    .X(_07821_));
 sky130_fd_sc_hd__mux4_2 _19539_ (.A0(\w[32][23] ),
    .A1(\w[36][23] ),
    .A2(\w[34][23] ),
    .A3(\w[38][23] ),
    .S0(net482),
    .S1(net488),
    .X(_07822_));
 sky130_fd_sc_hd__mux4_2 _19540_ (.A0(\w[40][23] ),
    .A1(\w[44][23] ),
    .A2(\w[42][23] ),
    .A3(\w[46][23] ),
    .S0(net482),
    .S1(net488),
    .X(_07823_));
 sky130_fd_sc_hd__mux4_2 _19541_ (.A0(\w[48][23] ),
    .A1(\w[52][23] ),
    .A2(\w[50][23] ),
    .A3(\w[54][23] ),
    .S0(net482),
    .S1(net488),
    .X(_07824_));
 sky130_fd_sc_hd__mux4_2 _19542_ (.A0(\w[56][23] ),
    .A1(\w[60][23] ),
    .A2(\w[58][23] ),
    .A3(\w[62][23] ),
    .S0(net482),
    .S1(net488),
    .X(_07825_));
 sky130_fd_sc_hd__mux4_2 _19543_ (.A0(_07822_),
    .A1(_07823_),
    .A2(_07824_),
    .A3(_07825_),
    .S0(net476),
    .S1(net474),
    .X(_07826_));
 sky130_fd_sc_hd__mux2i_4 _19544_ (.A0(_07821_),
    .A1(_07826_),
    .S(net473),
    .Y(_11765_));
 sky130_fd_sc_hd__mux4_2 _19545_ (.A0(\w[0][24] ),
    .A1(\w[4][24] ),
    .A2(\w[2][24] ),
    .A3(\w[6][24] ),
    .S0(net479),
    .S1(net489),
    .X(_07827_));
 sky130_fd_sc_hd__mux4_2 _19546_ (.A0(\w[8][24] ),
    .A1(\w[12][24] ),
    .A2(\w[10][24] ),
    .A3(\w[14][24] ),
    .S0(net479),
    .S1(net489),
    .X(_07828_));
 sky130_fd_sc_hd__mux4_2 _19547_ (.A0(\w[16][24] ),
    .A1(\w[20][24] ),
    .A2(\w[18][24] ),
    .A3(\w[22][24] ),
    .S0(net479),
    .S1(net489),
    .X(_07829_));
 sky130_fd_sc_hd__mux4_2 _19548_ (.A0(\w[24][24] ),
    .A1(\w[28][24] ),
    .A2(\w[26][24] ),
    .A3(\w[30][24] ),
    .S0(net479),
    .S1(net489),
    .X(_07830_));
 sky130_fd_sc_hd__mux4_2 _19549_ (.A0(_07827_),
    .A1(_07828_),
    .A2(_07829_),
    .A3(_07830_),
    .S0(net477),
    .S1(net475),
    .X(_07831_));
 sky130_fd_sc_hd__mux4_2 _19550_ (.A0(\w[32][24] ),
    .A1(\w[36][24] ),
    .A2(\w[34][24] ),
    .A3(\w[38][24] ),
    .S0(net480),
    .S1(net489),
    .X(_07832_));
 sky130_fd_sc_hd__mux4_2 _19551_ (.A0(\w[40][24] ),
    .A1(\w[44][24] ),
    .A2(\w[42][24] ),
    .A3(\w[46][24] ),
    .S0(net479),
    .S1(net489),
    .X(_07833_));
 sky130_fd_sc_hd__mux4_2 _19552_ (.A0(\w[48][24] ),
    .A1(\w[52][24] ),
    .A2(\w[50][24] ),
    .A3(\w[54][24] ),
    .S0(net480),
    .S1(net489),
    .X(_07834_));
 sky130_fd_sc_hd__mux4_2 _19553_ (.A0(\w[56][24] ),
    .A1(\w[60][24] ),
    .A2(\w[58][24] ),
    .A3(\w[62][24] ),
    .S0(net480),
    .S1(net489),
    .X(_07835_));
 sky130_fd_sc_hd__mux4_2 _19554_ (.A0(_07832_),
    .A1(_07833_),
    .A2(_07834_),
    .A3(_07835_),
    .S0(net477),
    .S1(net475),
    .X(_07836_));
 sky130_fd_sc_hd__mux2i_4 _19555_ (.A0(_07831_),
    .A1(_07836_),
    .S(net473),
    .Y(_11773_));
 sky130_fd_sc_hd__mux4_2 _19556_ (.A0(\w[0][25] ),
    .A1(\w[4][25] ),
    .A2(\w[2][25] ),
    .A3(\w[6][25] ),
    .S0(net482),
    .S1(net487),
    .X(_07837_));
 sky130_fd_sc_hd__mux4_2 _19557_ (.A0(\w[8][25] ),
    .A1(\w[12][25] ),
    .A2(\w[10][25] ),
    .A3(\w[14][25] ),
    .S0(net482),
    .S1(net487),
    .X(_07838_));
 sky130_fd_sc_hd__mux4_2 _19558_ (.A0(\w[16][25] ),
    .A1(\w[20][25] ),
    .A2(\w[18][25] ),
    .A3(\w[22][25] ),
    .S0(net481),
    .S1(net487),
    .X(_07839_));
 sky130_fd_sc_hd__mux4_2 _19559_ (.A0(\w[24][25] ),
    .A1(\w[28][25] ),
    .A2(\w[26][25] ),
    .A3(\w[30][25] ),
    .S0(net481),
    .S1(net487),
    .X(_07840_));
 sky130_fd_sc_hd__mux4_2 _19560_ (.A0(_07837_),
    .A1(_07838_),
    .A2(_07839_),
    .A3(_07840_),
    .S0(net476),
    .S1(net475),
    .X(_07841_));
 sky130_fd_sc_hd__mux4_2 _19561_ (.A0(\w[32][25] ),
    .A1(\w[36][25] ),
    .A2(\w[34][25] ),
    .A3(\w[38][25] ),
    .S0(net481),
    .S1(net488),
    .X(_07842_));
 sky130_fd_sc_hd__mux4_2 _19562_ (.A0(\w[40][25] ),
    .A1(\w[44][25] ),
    .A2(\w[42][25] ),
    .A3(\w[46][25] ),
    .S0(net481),
    .S1(net488),
    .X(_07843_));
 sky130_fd_sc_hd__mux4_2 _19563_ (.A0(\w[48][25] ),
    .A1(\w[52][25] ),
    .A2(\w[50][25] ),
    .A3(\w[54][25] ),
    .S0(net481),
    .S1(net488),
    .X(_07844_));
 sky130_fd_sc_hd__mux4_2 _19564_ (.A0(\w[56][25] ),
    .A1(\w[60][25] ),
    .A2(\w[58][25] ),
    .A3(\w[62][25] ),
    .S0(net481),
    .S1(net488),
    .X(_07845_));
 sky130_fd_sc_hd__mux4_2 _19565_ (.A0(_07842_),
    .A1(_07843_),
    .A2(_07844_),
    .A3(_07845_),
    .S0(net476),
    .S1(net475),
    .X(_07846_));
 sky130_fd_sc_hd__mux2i_4 _19566_ (.A0(_07841_),
    .A1(_07846_),
    .S(net473),
    .Y(_11781_));
 sky130_fd_sc_hd__mux4_2 _19567_ (.A0(\w[0][26] ),
    .A1(\w[4][26] ),
    .A2(\w[2][26] ),
    .A3(\w[6][26] ),
    .S0(net482),
    .S1(net487),
    .X(_07847_));
 sky130_fd_sc_hd__mux4_2 _19568_ (.A0(\w[8][26] ),
    .A1(\w[12][26] ),
    .A2(\w[10][26] ),
    .A3(\w[14][26] ),
    .S0(net482),
    .S1(net487),
    .X(_07848_));
 sky130_fd_sc_hd__mux4_2 _19569_ (.A0(\w[16][26] ),
    .A1(\w[20][26] ),
    .A2(\w[18][26] ),
    .A3(\w[22][26] ),
    .S0(net482),
    .S1(net487),
    .X(_07849_));
 sky130_fd_sc_hd__mux4_2 _19570_ (.A0(\w[24][26] ),
    .A1(\w[28][26] ),
    .A2(\w[26][26] ),
    .A3(\w[30][26] ),
    .S0(net482),
    .S1(net487),
    .X(_07850_));
 sky130_fd_sc_hd__mux4_2 _19571_ (.A0(_07847_),
    .A1(_07848_),
    .A2(_07849_),
    .A3(_07850_),
    .S0(net476),
    .S1(net475),
    .X(_07851_));
 sky130_fd_sc_hd__mux4_2 _19572_ (.A0(\w[32][26] ),
    .A1(\w[36][26] ),
    .A2(\w[34][26] ),
    .A3(\w[38][26] ),
    .S0(net481),
    .S1(net488),
    .X(_07852_));
 sky130_fd_sc_hd__mux4_2 _19573_ (.A0(\w[40][26] ),
    .A1(\w[44][26] ),
    .A2(\w[42][26] ),
    .A3(\w[46][26] ),
    .S0(net481),
    .S1(net488),
    .X(_07853_));
 sky130_fd_sc_hd__mux4_2 _19574_ (.A0(\w[48][26] ),
    .A1(\w[52][26] ),
    .A2(\w[50][26] ),
    .A3(\w[54][26] ),
    .S0(net481),
    .S1(net488),
    .X(_07854_));
 sky130_fd_sc_hd__mux4_2 _19575_ (.A0(\w[56][26] ),
    .A1(\w[60][26] ),
    .A2(\w[58][26] ),
    .A3(\w[62][26] ),
    .S0(net481),
    .S1(net488),
    .X(_07855_));
 sky130_fd_sc_hd__mux4_2 _19576_ (.A0(_07852_),
    .A1(_07853_),
    .A2(_07854_),
    .A3(_07855_),
    .S0(net476),
    .S1(net475),
    .X(_07856_));
 sky130_fd_sc_hd__mux2i_4 _19577_ (.A0(_07851_),
    .A1(_07856_),
    .S(net473),
    .Y(_11789_));
 sky130_fd_sc_hd__mux4_2 _19578_ (.A0(\w[0][27] ),
    .A1(\w[4][27] ),
    .A2(\w[2][27] ),
    .A3(\w[6][27] ),
    .S0(net483),
    .S1(net491),
    .X(_07857_));
 sky130_fd_sc_hd__mux4_2 _19579_ (.A0(\w[8][27] ),
    .A1(\w[12][27] ),
    .A2(\w[10][27] ),
    .A3(\w[14][27] ),
    .S0(net483),
    .S1(net491),
    .X(_07858_));
 sky130_fd_sc_hd__mux4_2 _19580_ (.A0(\w[16][27] ),
    .A1(\w[20][27] ),
    .A2(\w[18][27] ),
    .A3(\w[22][27] ),
    .S0(net483),
    .S1(net491),
    .X(_07859_));
 sky130_fd_sc_hd__mux4_2 _19581_ (.A0(\w[24][27] ),
    .A1(\w[28][27] ),
    .A2(\w[26][27] ),
    .A3(\w[30][27] ),
    .S0(net483),
    .S1(net491),
    .X(_07860_));
 sky130_fd_sc_hd__mux4_2 _19582_ (.A0(_07857_),
    .A1(_07858_),
    .A2(_07859_),
    .A3(_07860_),
    .S0(net476),
    .S1(net474),
    .X(_07861_));
 sky130_fd_sc_hd__mux4_2 _19583_ (.A0(\w[32][27] ),
    .A1(\w[36][27] ),
    .A2(\w[34][27] ),
    .A3(\w[38][27] ),
    .S0(net483),
    .S1(net491),
    .X(_07862_));
 sky130_fd_sc_hd__mux4_2 _19584_ (.A0(\w[40][27] ),
    .A1(\w[44][27] ),
    .A2(\w[42][27] ),
    .A3(\w[46][27] ),
    .S0(net483),
    .S1(net491),
    .X(_07863_));
 sky130_fd_sc_hd__mux4_2 _19585_ (.A0(\w[48][27] ),
    .A1(\w[52][27] ),
    .A2(\w[50][27] ),
    .A3(\w[54][27] ),
    .S0(net483),
    .S1(net491),
    .X(_07864_));
 sky130_fd_sc_hd__mux4_2 _19586_ (.A0(\w[56][27] ),
    .A1(\w[60][27] ),
    .A2(\w[58][27] ),
    .A3(\w[62][27] ),
    .S0(net483),
    .S1(net491),
    .X(_07865_));
 sky130_fd_sc_hd__mux4_2 _19587_ (.A0(_07862_),
    .A1(_07863_),
    .A2(_07864_),
    .A3(_07865_),
    .S0(net476),
    .S1(net474),
    .X(_07866_));
 sky130_fd_sc_hd__mux2i_4 _19588_ (.A0(_07861_),
    .A1(_07866_),
    .S(net473),
    .Y(_11797_));
 sky130_fd_sc_hd__mux4_2 _19589_ (.A0(\w[0][28] ),
    .A1(\w[4][28] ),
    .A2(\w[2][28] ),
    .A3(\w[6][28] ),
    .S0(net483),
    .S1(net491),
    .X(_07867_));
 sky130_fd_sc_hd__mux4_2 _19590_ (.A0(\w[8][28] ),
    .A1(\w[12][28] ),
    .A2(\w[10][28] ),
    .A3(\w[14][28] ),
    .S0(net483),
    .S1(net491),
    .X(_07868_));
 sky130_fd_sc_hd__mux4_2 _19591_ (.A0(\w[16][28] ),
    .A1(\w[20][28] ),
    .A2(\w[18][28] ),
    .A3(\w[22][28] ),
    .S0(net483),
    .S1(net491),
    .X(_07869_));
 sky130_fd_sc_hd__mux4_2 _19592_ (.A0(\w[24][28] ),
    .A1(\w[28][28] ),
    .A2(\w[26][28] ),
    .A3(\w[30][28] ),
    .S0(net483),
    .S1(net491),
    .X(_07870_));
 sky130_fd_sc_hd__mux4_2 _19593_ (.A0(_07867_),
    .A1(_07868_),
    .A2(_07869_),
    .A3(_07870_),
    .S0(net476),
    .S1(net474),
    .X(_07871_));
 sky130_fd_sc_hd__mux4_2 _19594_ (.A0(\w[32][28] ),
    .A1(\w[36][28] ),
    .A2(\w[34][28] ),
    .A3(\w[38][28] ),
    .S0(net482),
    .S1(net488),
    .X(_07872_));
 sky130_fd_sc_hd__mux4_2 _19595_ (.A0(\w[40][28] ),
    .A1(\w[44][28] ),
    .A2(\w[42][28] ),
    .A3(\w[46][28] ),
    .S0(net482),
    .S1(net487),
    .X(_07873_));
 sky130_fd_sc_hd__mux4_2 _19596_ (.A0(\w[48][28] ),
    .A1(\w[52][28] ),
    .A2(\w[50][28] ),
    .A3(\w[54][28] ),
    .S0(net482),
    .S1(net487),
    .X(_07874_));
 sky130_fd_sc_hd__mux4_2 _19597_ (.A0(\w[56][28] ),
    .A1(\w[60][28] ),
    .A2(\w[58][28] ),
    .A3(\w[62][28] ),
    .S0(net482),
    .S1(net488),
    .X(_07875_));
 sky130_fd_sc_hd__mux4_2 _19598_ (.A0(_07872_),
    .A1(_07873_),
    .A2(_07874_),
    .A3(_07875_),
    .S0(net476),
    .S1(net474),
    .X(_07876_));
 sky130_fd_sc_hd__mux2i_4 _19599_ (.A0(_07871_),
    .A1(_07876_),
    .S(net473),
    .Y(_11805_));
 sky130_fd_sc_hd__mux4_2 _19600_ (.A0(\w[0][29] ),
    .A1(\w[4][29] ),
    .A2(\w[2][29] ),
    .A3(\w[6][29] ),
    .S0(net478),
    .S1(net486),
    .X(_07877_));
 sky130_fd_sc_hd__mux4_2 _19601_ (.A0(\w[8][29] ),
    .A1(\w[12][29] ),
    .A2(\w[10][29] ),
    .A3(\w[14][29] ),
    .S0(net478),
    .S1(net486),
    .X(_07878_));
 sky130_fd_sc_hd__mux4_2 _19602_ (.A0(\w[16][29] ),
    .A1(\w[20][29] ),
    .A2(\w[18][29] ),
    .A3(\w[22][29] ),
    .S0(net478),
    .S1(net486),
    .X(_07879_));
 sky130_fd_sc_hd__mux4_2 _19603_ (.A0(\w[24][29] ),
    .A1(\w[28][29] ),
    .A2(\w[26][29] ),
    .A3(\w[30][29] ),
    .S0(net478),
    .S1(net486),
    .X(_07880_));
 sky130_fd_sc_hd__mux4_2 _19604_ (.A0(_07877_),
    .A1(_07878_),
    .A2(_07879_),
    .A3(_07880_),
    .S0(net546),
    .S1(net474),
    .X(_07881_));
 sky130_fd_sc_hd__mux4_2 _19605_ (.A0(\w[32][29] ),
    .A1(\w[36][29] ),
    .A2(\w[34][29] ),
    .A3(\w[38][29] ),
    .S0(net478),
    .S1(net486),
    .X(_07882_));
 sky130_fd_sc_hd__mux4_2 _19606_ (.A0(\w[40][29] ),
    .A1(\w[44][29] ),
    .A2(\w[42][29] ),
    .A3(\w[46][29] ),
    .S0(net478),
    .S1(net486),
    .X(_07883_));
 sky130_fd_sc_hd__mux4_2 _19607_ (.A0(\w[48][29] ),
    .A1(\w[52][29] ),
    .A2(\w[50][29] ),
    .A3(\w[54][29] ),
    .S0(net478),
    .S1(net486),
    .X(_07884_));
 sky130_fd_sc_hd__mux4_2 _19608_ (.A0(\w[56][29] ),
    .A1(\w[60][29] ),
    .A2(\w[58][29] ),
    .A3(\w[62][29] ),
    .S0(net478),
    .S1(net486),
    .X(_07885_));
 sky130_fd_sc_hd__mux4_2 _19609_ (.A0(_07882_),
    .A1(_07883_),
    .A2(_07884_),
    .A3(_07885_),
    .S0(net546),
    .S1(net474),
    .X(_07886_));
 sky130_fd_sc_hd__mux2i_4 _19610_ (.A0(_07881_),
    .A1(_07886_),
    .S(net545),
    .Y(_11813_));
 sky130_fd_sc_hd__mux4_2 _19611_ (.A0(\w[0][30] ),
    .A1(\w[4][30] ),
    .A2(\w[2][30] ),
    .A3(\w[6][30] ),
    .S0(net478),
    .S1(net486),
    .X(_07887_));
 sky130_fd_sc_hd__mux4_2 _19612_ (.A0(\w[8][30] ),
    .A1(\w[12][30] ),
    .A2(\w[10][30] ),
    .A3(\w[14][30] ),
    .S0(net478),
    .S1(net486),
    .X(_07888_));
 sky130_fd_sc_hd__mux4_2 _19613_ (.A0(\w[16][30] ),
    .A1(\w[20][30] ),
    .A2(\w[18][30] ),
    .A3(\w[22][30] ),
    .S0(net478),
    .S1(net486),
    .X(_07889_));
 sky130_fd_sc_hd__mux4_2 _19614_ (.A0(\w[24][30] ),
    .A1(\w[28][30] ),
    .A2(\w[26][30] ),
    .A3(\w[30][30] ),
    .S0(net478),
    .S1(net486),
    .X(_07890_));
 sky130_fd_sc_hd__mux4_2 _19615_ (.A0(_07887_),
    .A1(_07888_),
    .A2(_07889_),
    .A3(_07890_),
    .S0(net546),
    .S1(net474),
    .X(_07891_));
 sky130_fd_sc_hd__mux4_2 _19616_ (.A0(\w[32][30] ),
    .A1(\w[36][30] ),
    .A2(\w[34][30] ),
    .A3(\w[38][30] ),
    .S0(net478),
    .S1(net486),
    .X(_07892_));
 sky130_fd_sc_hd__mux4_2 _19617_ (.A0(\w[40][30] ),
    .A1(\w[44][30] ),
    .A2(\w[42][30] ),
    .A3(\w[46][30] ),
    .S0(net478),
    .S1(net486),
    .X(_07893_));
 sky130_fd_sc_hd__mux4_2 _19618_ (.A0(\w[48][30] ),
    .A1(\w[52][30] ),
    .A2(\w[50][30] ),
    .A3(\w[54][30] ),
    .S0(net478),
    .S1(net486),
    .X(_07894_));
 sky130_fd_sc_hd__mux4_2 _19619_ (.A0(\w[56][30] ),
    .A1(\w[60][30] ),
    .A2(\w[58][30] ),
    .A3(\w[62][30] ),
    .S0(net478),
    .S1(net486),
    .X(_07895_));
 sky130_fd_sc_hd__mux4_2 _19620_ (.A0(_07892_),
    .A1(_07893_),
    .A2(_07894_),
    .A3(_07895_),
    .S0(net546),
    .S1(net474),
    .X(_07896_));
 sky130_fd_sc_hd__mux2i_4 _19621_ (.A0(_07891_),
    .A1(_07896_),
    .S(net545),
    .Y(_11821_));
 sky130_fd_sc_hd__inv_1 _19622_ (.A(_12504_),
    .Y(_12662_));
 sky130_fd_sc_hd__inv_1 _19623_ (.A(_12883_),
    .Y(\hash.CA1.p1[1] ));
 sky130_fd_sc_hd__inv_1 _19624_ (.A(_12886_),
    .Y(\hash.CA1.p2[2] ));
 sky130_fd_sc_hd__inv_1 _19625_ (.A(_12893_),
    .Y(\hash.CA1.p3[2] ));
 sky130_fd_sc_hd__inv_1 _19626_ (.A(_12897_),
    .Y(\hash.CA1.p5[1] ));
 sky130_fd_sc_hd__inv_1 _19627_ (.A(_12104_),
    .Y(_12107_));
 sky130_fd_sc_hd__inv_1 _19628_ (.A(_12512_),
    .Y(_12891_));
 sky130_fd_sc_hd__inv_1 _19629_ (.A(_12659_),
    .Y(_12661_));
 sky130_fd_sc_hd__inv_1 _19630_ (.A(_12686_),
    .Y(_12687_));
 sky130_fd_sc_hd__inv_1 _19631_ (.A(_12874_),
    .Y(_12876_));
 sky130_fd_sc_hd__inv_1 _19632_ (.A(_12094_),
    .Y(_12106_));
 sky130_fd_sc_hd__inv_1 _19633_ (.A(_12506_),
    .Y(_12890_));
 sky130_fd_sc_hd__inv_1 _19634_ (.A(_12655_),
    .Y(_12660_));
 sky130_fd_sc_hd__inv_1 _19635_ (.A(_12658_),
    .Y(_12670_));
 sky130_fd_sc_hd__inv_1 _19636_ (.A(_12685_),
    .Y(_12696_));
 sky130_fd_sc_hd__inv_1 _19637_ (.A(_12865_),
    .Y(_12875_));
 sky130_fd_sc_hd__clkinvlp_4 _19638_ (.A(\count_hash2[1] ),
    .Y(_00656_));
 sky130_fd_sc_hd__inv_6 _19639_ (.A(net371),
    .Y(_00654_));
 sky130_fd_sc_hd__xor2_1 _19640_ (.A(_11335_),
    .B(_02699_),
    .X(_07897_));
 sky130_fd_sc_hd__xnor2_1 _19641_ (.A(_11090_),
    .B(_07897_),
    .Y(_12983_));
 sky130_fd_sc_hd__inv_1 _19642_ (.A(_11590_),
    .Y(_12990_));
 sky130_fd_sc_hd__inv_1 _19643_ (.A(_11598_),
    .Y(_12994_));
 sky130_fd_sc_hd__inv_1 _19644_ (.A(_11609_),
    .Y(_12998_));
 sky130_fd_sc_hd__inv_1 _19645_ (.A(_11617_),
    .Y(_13002_));
 sky130_fd_sc_hd__inv_1 _19646_ (.A(_11625_),
    .Y(_13006_));
 sky130_fd_sc_hd__clkinv_2 _19647_ (.A(_11633_),
    .Y(_13010_));
 sky130_fd_sc_hd__inv_2 _19648_ (.A(_11641_),
    .Y(_13014_));
 sky130_fd_sc_hd__clkinv_1 _19649_ (.A(_11649_),
    .Y(_13018_));
 sky130_fd_sc_hd__clkinv_1 _19650_ (.A(_11657_),
    .Y(_13022_));
 sky130_fd_sc_hd__clkinv_1 _19651_ (.A(_11665_),
    .Y(_13026_));
 sky130_fd_sc_hd__inv_1 _19652_ (.A(_11673_),
    .Y(_13030_));
 sky130_fd_sc_hd__inv_1 _19653_ (.A(_11681_),
    .Y(_13034_));
 sky130_fd_sc_hd__inv_1 _19654_ (.A(_11689_),
    .Y(_13038_));
 sky130_fd_sc_hd__inv_1 _19655_ (.A(_11697_),
    .Y(_13042_));
 sky130_fd_sc_hd__inv_1 _19656_ (.A(_11705_),
    .Y(_13046_));
 sky130_fd_sc_hd__inv_1 _19657_ (.A(_11713_),
    .Y(_13050_));
 sky130_fd_sc_hd__inv_1 _19658_ (.A(_11721_),
    .Y(_13054_));
 sky130_fd_sc_hd__inv_1 _19659_ (.A(_11729_),
    .Y(_13058_));
 sky130_fd_sc_hd__clkinv_1 _19660_ (.A(_11737_),
    .Y(_13062_));
 sky130_fd_sc_hd__inv_1 _19661_ (.A(_11745_),
    .Y(_13066_));
 sky130_fd_sc_hd__clkinv_1 _19662_ (.A(_11753_),
    .Y(_13070_));
 sky130_fd_sc_hd__inv_1 _19663_ (.A(_11761_),
    .Y(_13074_));
 sky130_fd_sc_hd__inv_1 _19664_ (.A(_11769_),
    .Y(_13078_));
 sky130_fd_sc_hd__inv_1 _19665_ (.A(_11777_),
    .Y(_13082_));
 sky130_fd_sc_hd__clkinv_1 _19666_ (.A(_11785_),
    .Y(_13086_));
 sky130_fd_sc_hd__clkinv_1 _19667_ (.A(_11793_),
    .Y(_13090_));
 sky130_fd_sc_hd__clkinv_1 _19668_ (.A(_11801_),
    .Y(_13094_));
 sky130_fd_sc_hd__clkinv_1 _19669_ (.A(_11809_),
    .Y(_13098_));
 sky130_fd_sc_hd__clkinv_1 _19670_ (.A(_11817_),
    .Y(_13102_));
 sky130_fd_sc_hd__mux4_2 _19671_ (.A0(\w[1][0] ),
    .A1(\w[5][0] ),
    .A2(\w[3][0] ),
    .A3(\w[7][0] ),
    .S0(net460),
    .S1(net470),
    .X(_07898_));
 sky130_fd_sc_hd__mux4_2 _19672_ (.A0(\w[9][0] ),
    .A1(\w[13][0] ),
    .A2(\w[11][0] ),
    .A3(\w[15][0] ),
    .S0(net460),
    .S1(net470),
    .X(_07899_));
 sky130_fd_sc_hd__mux4_2 _19673_ (.A0(\w[17][0] ),
    .A1(\w[21][0] ),
    .A2(\w[19][0] ),
    .A3(\w[23][0] ),
    .S0(net460),
    .S1(net470),
    .X(_07900_));
 sky130_fd_sc_hd__mux4_2 _19674_ (.A0(\w[25][0] ),
    .A1(\w[29][0] ),
    .A2(\w[27][0] ),
    .A3(\w[31][0] ),
    .S0(net460),
    .S1(net470),
    .X(_07901_));
 sky130_fd_sc_hd__mux4_2 _19675_ (.A0(_07898_),
    .A1(_07899_),
    .A2(_07900_),
    .A3(_07901_),
    .S0(net456),
    .S1(net454),
    .X(_07902_));
 sky130_fd_sc_hd__mux4_2 _19676_ (.A0(\w[33][0] ),
    .A1(\w[37][0] ),
    .A2(\w[35][0] ),
    .A3(\w[39][0] ),
    .S0(net460),
    .S1(net469),
    .X(_07903_));
 sky130_fd_sc_hd__mux4_2 _19677_ (.A0(\w[41][0] ),
    .A1(\w[45][0] ),
    .A2(\w[43][0] ),
    .A3(\w[47][0] ),
    .S0(net460),
    .S1(net469),
    .X(_07904_));
 sky130_fd_sc_hd__mux4_2 _19678_ (.A0(\w[49][0] ),
    .A1(\w[53][0] ),
    .A2(\w[51][0] ),
    .A3(\w[55][0] ),
    .S0(net460),
    .S1(net469),
    .X(_07905_));
 sky130_fd_sc_hd__mux4_2 _19679_ (.A0(\w[57][0] ),
    .A1(\w[61][0] ),
    .A2(\w[59][0] ),
    .A3(\w[63][0] ),
    .S0(net460),
    .S1(net469),
    .X(_07906_));
 sky130_fd_sc_hd__mux4_2 _19680_ (.A0(_07903_),
    .A1(_07904_),
    .A2(_07905_),
    .A3(_07906_),
    .S0(net456),
    .S1(net454),
    .X(_07907_));
 sky130_fd_sc_hd__mux2_8 _19681_ (.A0(_07902_),
    .A1(_07907_),
    .S(net453),
    .X(_13106_));
 sky130_fd_sc_hd__inv_1 _19682_ (.A(_11838_),
    .Y(_13113_));
 sky130_fd_sc_hd__inv_1 _19683_ (.A(_11846_),
    .Y(_13117_));
 sky130_fd_sc_hd__inv_1 _19684_ (.A(_11857_),
    .Y(_13121_));
 sky130_fd_sc_hd__inv_1 _19685_ (.A(_11865_),
    .Y(_13125_));
 sky130_fd_sc_hd__inv_1 _19686_ (.A(_11873_),
    .Y(_13129_));
 sky130_fd_sc_hd__inv_1 _19687_ (.A(_11881_),
    .Y(_13133_));
 sky130_fd_sc_hd__clkinv_2 _19688_ (.A(_11889_),
    .Y(_13137_));
 sky130_fd_sc_hd__clkinv_1 _19689_ (.A(_11897_),
    .Y(_13141_));
 sky130_fd_sc_hd__inv_2 _19690_ (.A(_11905_),
    .Y(_13145_));
 sky130_fd_sc_hd__clkinv_1 _19691_ (.A(_11913_),
    .Y(_13149_));
 sky130_fd_sc_hd__inv_1 _19692_ (.A(_11921_),
    .Y(_13153_));
 sky130_fd_sc_hd__inv_1 _19693_ (.A(_11929_),
    .Y(_13157_));
 sky130_fd_sc_hd__inv_1 _19694_ (.A(_11937_),
    .Y(_13161_));
 sky130_fd_sc_hd__inv_1 _19695_ (.A(_11945_),
    .Y(_13165_));
 sky130_fd_sc_hd__inv_1 _19696_ (.A(_11953_),
    .Y(_13169_));
 sky130_fd_sc_hd__clkinv_1 _19697_ (.A(_11961_),
    .Y(_13173_));
 sky130_fd_sc_hd__clkinv_1 _19698_ (.A(_11969_),
    .Y(_13177_));
 sky130_fd_sc_hd__clkinv_1 _19699_ (.A(_11977_),
    .Y(_13181_));
 sky130_fd_sc_hd__inv_1 _19700_ (.A(_11985_),
    .Y(_13185_));
 sky130_fd_sc_hd__inv_1 _19701_ (.A(_11993_),
    .Y(_13189_));
 sky130_fd_sc_hd__clkinv_1 _19702_ (.A(_12001_),
    .Y(_13193_));
 sky130_fd_sc_hd__clkinv_1 _19703_ (.A(_12009_),
    .Y(_13197_));
 sky130_fd_sc_hd__inv_1 _19704_ (.A(_12017_),
    .Y(_13201_));
 sky130_fd_sc_hd__inv_1 _19705_ (.A(_12025_),
    .Y(_13205_));
 sky130_fd_sc_hd__inv_2 _19706_ (.A(_12033_),
    .Y(_13209_));
 sky130_fd_sc_hd__clkinv_1 _19707_ (.A(_12041_),
    .Y(_13213_));
 sky130_fd_sc_hd__inv_1 _19708_ (.A(_12049_),
    .Y(_13217_));
 sky130_fd_sc_hd__inv_1 _19709_ (.A(_12057_),
    .Y(_13221_));
 sky130_fd_sc_hd__inv_1 _19710_ (.A(_12065_),
    .Y(_13225_));
 sky130_fd_sc_hd__mux2_4 _19711_ (.A0(\hash.CA2.f_dash[0] ),
    .A1(\hash.CA2.e_dash[0] ),
    .S(\hash.CA2.S1.X[0] ),
    .X(_13229_));
 sky130_fd_sc_hd__inv_1 _19712_ (.A(_12078_),
    .Y(_12092_));
 sky130_fd_sc_hd__mux2_4 _19713_ (.A0(\hash.CA2.f_dash[2] ),
    .A1(\hash.CA2.e_dash[2] ),
    .S(\hash.CA2.S1.X[2] ),
    .X(_13242_));
 sky130_fd_sc_hd__inv_1 _19714_ (.A(_12090_),
    .Y(_12101_));
 sky130_fd_sc_hd__mux2_1 _19715_ (.A0(\hash.CA2.f_dash[3] ),
    .A1(\hash.CA2.e_dash[3] ),
    .S(\hash.CA2.S1.X[3] ),
    .X(_13249_));
 sky130_fd_sc_hd__inv_1 _19716_ (.A(_12099_),
    .Y(_12115_));
 sky130_fd_sc_hd__mux2_1 _19717_ (.A0(\hash.CA2.f_dash[4] ),
    .A1(\hash.CA2.e_dash[4] ),
    .S(\hash.CA2.S1.X[4] ),
    .X(_13256_));
 sky130_fd_sc_hd__inv_2 _19718_ (.A(_12113_),
    .Y(_12124_));
 sky130_fd_sc_hd__mux2_4 _19719_ (.A0(\hash.CA2.f_dash[5] ),
    .A1(\hash.CA2.e_dash[5] ),
    .S(\hash.CA2.S1.X[5] ),
    .X(_13263_));
 sky130_fd_sc_hd__inv_1 _19720_ (.A(_12122_),
    .Y(_12133_));
 sky130_fd_sc_hd__mux2_8 _19721_ (.A0(\hash.CA2.f_dash[6] ),
    .A1(\hash.CA2.e_dash[6] ),
    .S(net1075),
    .X(_13270_));
 sky130_fd_sc_hd__inv_1 _19722_ (.A(_12131_),
    .Y(_12142_));
 sky130_fd_sc_hd__mux2_8 _19723_ (.A0(\hash.CA2.f_dash[7] ),
    .A1(\hash.CA2.e_dash[7] ),
    .S(net1081),
    .X(_13277_));
 sky130_fd_sc_hd__inv_1 _19724_ (.A(_12140_),
    .Y(_12151_));
 sky130_fd_sc_hd__mux2_8 _19725_ (.A0(\hash.CA2.f_dash[8] ),
    .A1(\hash.CA2.e_dash[8] ),
    .S(net1110),
    .X(_13284_));
 sky130_fd_sc_hd__inv_1 _19726_ (.A(_12149_),
    .Y(_12160_));
 sky130_fd_sc_hd__mux2_8 _19727_ (.A0(\hash.CA2.f_dash[9] ),
    .A1(\hash.CA2.e_dash[9] ),
    .S(\hash.CA2.S1.X[9] ),
    .X(_13291_));
 sky130_fd_sc_hd__inv_1 _19728_ (.A(_12158_),
    .Y(_12169_));
 sky130_fd_sc_hd__mux2_8 _19729_ (.A0(\hash.CA2.f_dash[10] ),
    .A1(\hash.CA2.e_dash[10] ),
    .S(\hash.CA2.S1.X[10] ),
    .X(_13298_));
 sky130_fd_sc_hd__inv_1 _19730_ (.A(_12167_),
    .Y(_12178_));
 sky130_fd_sc_hd__mux2_4 _19731_ (.A0(\hash.CA2.f_dash[11] ),
    .A1(\hash.CA2.e_dash[11] ),
    .S(\hash.CA2.S1.X[11] ),
    .X(_13305_));
 sky130_fd_sc_hd__inv_1 _19732_ (.A(_12176_),
    .Y(_12187_));
 sky130_fd_sc_hd__mux2_8 _19733_ (.A0(\hash.CA2.f_dash[12] ),
    .A1(\hash.CA2.e_dash[12] ),
    .S(\hash.CA2.S1.X[12] ),
    .X(_13312_));
 sky130_fd_sc_hd__inv_2 _19734_ (.A(_12185_),
    .Y(_12196_));
 sky130_fd_sc_hd__nand2_2 _19735_ (.A(\hash.CA2.S1.X[13] ),
    .B(\hash.CA2.e_dash[13] ),
    .Y(_07908_));
 sky130_fd_sc_hd__o21ai_4 _19736_ (.A1(\hash.CA2.S1.X[13] ),
    .A2(_06314_),
    .B1(_07908_),
    .Y(_13319_));
 sky130_fd_sc_hd__inv_1 _19737_ (.A(_12194_),
    .Y(_12205_));
 sky130_fd_sc_hd__mux2_8 _19738_ (.A0(\hash.CA2.f_dash[14] ),
    .A1(\hash.CA2.e_dash[14] ),
    .S(\hash.CA2.S1.X[14] ),
    .X(_13326_));
 sky130_fd_sc_hd__inv_1 _19739_ (.A(_12203_),
    .Y(_12214_));
 sky130_fd_sc_hd__mux2_8 _19740_ (.A0(\hash.CA2.f_dash[15] ),
    .A1(\hash.CA2.e_dash[15] ),
    .S(\hash.CA2.S1.X[15] ),
    .X(_13333_));
 sky130_fd_sc_hd__inv_1 _19741_ (.A(_12212_),
    .Y(_12223_));
 sky130_fd_sc_hd__mux2_8 _19742_ (.A0(\hash.CA2.f_dash[16] ),
    .A1(\hash.CA2.e_dash[16] ),
    .S(\hash.CA2.S1.X[16] ),
    .X(_13340_));
 sky130_fd_sc_hd__inv_1 _19743_ (.A(_12221_),
    .Y(_12232_));
 sky130_fd_sc_hd__mux2_8 _19744_ (.A0(\hash.CA2.f_dash[17] ),
    .A1(\hash.CA2.e_dash[17] ),
    .S(\hash.CA2.S1.X[17] ),
    .X(_13347_));
 sky130_fd_sc_hd__inv_1 _19745_ (.A(_12230_),
    .Y(_12241_));
 sky130_fd_sc_hd__mux2_8 _19746_ (.A0(\hash.CA2.f_dash[18] ),
    .A1(\hash.CA2.e_dash[18] ),
    .S(\hash.CA2.S1.X[18] ),
    .X(_13354_));
 sky130_fd_sc_hd__inv_1 _19747_ (.A(_12239_),
    .Y(_12250_));
 sky130_fd_sc_hd__mux2_8 _19748_ (.A0(\hash.CA2.f_dash[19] ),
    .A1(\hash.CA2.e_dash[19] ),
    .S(\hash.CA2.S1.X[19] ),
    .X(_13361_));
 sky130_fd_sc_hd__inv_1 _19749_ (.A(_12248_),
    .Y(_12259_));
 sky130_fd_sc_hd__mux2_8 _19750_ (.A0(\hash.CA2.f_dash[20] ),
    .A1(\hash.CA2.e_dash[20] ),
    .S(\hash.CA2.S1.X[20] ),
    .X(_13368_));
 sky130_fd_sc_hd__inv_1 _19751_ (.A(_12257_),
    .Y(_12268_));
 sky130_fd_sc_hd__mux2_8 _19752_ (.A0(\hash.CA2.f_dash[21] ),
    .A1(\hash.CA2.e_dash[21] ),
    .S(\hash.CA2.S1.X[21] ),
    .X(_13375_));
 sky130_fd_sc_hd__inv_1 _19753_ (.A(_12266_),
    .Y(_12277_));
 sky130_fd_sc_hd__mux2_8 _19754_ (.A0(\hash.CA2.f_dash[22] ),
    .A1(\hash.CA2.e_dash[22] ),
    .S(\hash.CA2.S1.X[22] ),
    .X(_13382_));
 sky130_fd_sc_hd__inv_1 _19755_ (.A(_12275_),
    .Y(_12286_));
 sky130_fd_sc_hd__mux2_8 _19756_ (.A0(\hash.CA2.f_dash[23] ),
    .A1(\hash.CA2.e_dash[23] ),
    .S(\hash.CA2.S1.X[23] ),
    .X(_13389_));
 sky130_fd_sc_hd__inv_1 _19757_ (.A(_12284_),
    .Y(_12295_));
 sky130_fd_sc_hd__mux2_8 _19758_ (.A0(\hash.CA2.f_dash[24] ),
    .A1(\hash.CA2.e_dash[24] ),
    .S(\hash.CA2.S1.X[24] ),
    .X(_13396_));
 sky130_fd_sc_hd__inv_1 _19759_ (.A(_12293_),
    .Y(_12304_));
 sky130_fd_sc_hd__mux2_8 _19760_ (.A0(\hash.CA2.f_dash[25] ),
    .A1(\hash.CA2.e_dash[25] ),
    .S(net1092),
    .X(_13403_));
 sky130_fd_sc_hd__inv_1 _19761_ (.A(_12302_),
    .Y(_12313_));
 sky130_fd_sc_hd__mux2_8 _19762_ (.A0(\hash.CA2.f_dash[26] ),
    .A1(\hash.CA2.e_dash[26] ),
    .S(net1100),
    .X(_13410_));
 sky130_fd_sc_hd__inv_1 _19763_ (.A(_12311_),
    .Y(_12322_));
 sky130_fd_sc_hd__mux2_8 _19764_ (.A0(\hash.CA2.f_dash[27] ),
    .A1(\hash.CA2.e_dash[27] ),
    .S(\hash.CA2.S1.X[27] ),
    .X(_13417_));
 sky130_fd_sc_hd__inv_1 _19765_ (.A(_12320_),
    .Y(_12331_));
 sky130_fd_sc_hd__mux2_8 _19766_ (.A0(\hash.CA2.f_dash[28] ),
    .A1(\hash.CA2.e_dash[28] ),
    .S(\hash.CA2.S1.X[28] ),
    .X(_13424_));
 sky130_fd_sc_hd__inv_1 _19767_ (.A(_12329_),
    .Y(_12340_));
 sky130_fd_sc_hd__mux2_4 _19768_ (.A0(\hash.CA2.f_dash[29] ),
    .A1(\hash.CA2.e_dash[29] ),
    .S(\hash.CA2.S1.X[29] ),
    .X(_13431_));
 sky130_fd_sc_hd__inv_1 _19769_ (.A(_12338_),
    .Y(_12349_));
 sky130_fd_sc_hd__mux2_8 _19770_ (.A0(\hash.CA2.f_dash[30] ),
    .A1(\hash.CA2.e_dash[30] ),
    .S(\hash.CA2.S1.X[30] ),
    .X(_13438_));
 sky130_fd_sc_hd__inv_1 _19771_ (.A(_12347_),
    .Y(_12358_));
 sky130_fd_sc_hd__inv_4 _19772_ (.A(\count_1[1] ),
    .Y(_00650_));
 sky130_fd_sc_hd__inv_4 _19773_ (.A(\count_2[1] ),
    .Y(_00652_));
 sky130_fd_sc_hd__a21oi_1 _19774_ (.A1(\hash.CA2.a_dash[2] ),
    .A2(_05998_),
    .B1(_04421_),
    .Y(_07909_));
 sky130_fd_sc_hd__nor2_1 _19775_ (.A(\hash.CA2.a_dash[2] ),
    .B(_05998_),
    .Y(_07910_));
 sky130_fd_sc_hd__o21ai_0 _19776_ (.A1(_07909_),
    .A2(_07910_),
    .B1(_06002_),
    .Y(_13551_));
 sky130_fd_sc_hd__o21ai_0 _19777_ (.A1(\hash.CA1.S0.X[3] ),
    .A2(\hash.CA1.b[3] ),
    .B1(\hash.CA2.a_dash[3] ),
    .Y(_07911_));
 sky130_fd_sc_hd__nand2_1 _19778_ (.A(_04470_),
    .B(\hash.CA1.S0.X[3] ),
    .Y(_07912_));
 sky130_fd_sc_hd__nand2_2 _19779_ (.A(_07911_),
    .B(_07912_),
    .Y(_13555_));
 sky130_fd_sc_hd__nor2_1 _19780_ (.A(_06010_),
    .B(\hash.CA1.b[4] ),
    .Y(_07913_));
 sky130_fd_sc_hd__a21oi_1 _19781_ (.A1(_04487_),
    .A2(_06010_),
    .B1(\hash.CA2.a_dash[4] ),
    .Y(_07914_));
 sky130_fd_sc_hd__nor2_1 _19782_ (.A(_07913_),
    .B(_07914_),
    .Y(_13559_));
 sky130_fd_sc_hd__nor2_1 _19783_ (.A(net340),
    .B(_04501_),
    .Y(_07915_));
 sky130_fd_sc_hd__nor2_1 _19784_ (.A(_06016_),
    .B(_07915_),
    .Y(_07916_));
 sky130_fd_sc_hd__o22a_1 _19785_ (.A1(\hash.CA1.S0.X[5] ),
    .A2(\hash.CA1.b[5] ),
    .B1(_07916_),
    .B2(\hash.CA2.a_dash[5] ),
    .X(_13563_));
 sky130_fd_sc_hd__nor2_1 _19786_ (.A(net340),
    .B(_04522_),
    .Y(_07917_));
 sky130_fd_sc_hd__o21ai_0 _19787_ (.A1(\hash.CA1.S0.X[6] ),
    .A2(\hash.CA1.b[6] ),
    .B1(\hash.CA2.a_dash[6] ),
    .Y(_07918_));
 sky130_fd_sc_hd__o21ai_0 _19788_ (.A1(_06024_),
    .A2(_07917_),
    .B1(_07918_),
    .Y(_13567_));
 sky130_fd_sc_hd__nand2_2 _19789_ (.A(_06030_),
    .B(_06031_),
    .Y(_07919_));
 sky130_fd_sc_hd__a21oi_1 _19790_ (.A1(\hash.CA1.S0.X[7] ),
    .A2(\hash.CA1.b[7] ),
    .B1(\hash.CA2.a_dash[7] ),
    .Y(_07920_));
 sky130_fd_sc_hd__a211oi_1 _19791_ (.A1(_04543_),
    .A2(_07919_),
    .B1(_07920_),
    .C1(net340),
    .Y(_13571_));
 sky130_fd_sc_hd__maj3_1 _19792_ (.A(\hash.CA2.a_dash[8] ),
    .B(_06043_),
    .C(_06279_),
    .X(_13575_));
 sky130_fd_sc_hd__maj3_4 _19793_ (.A(\hash.CA2.a_dash[9] ),
    .B(\hash.CA1.S0.X[9] ),
    .C(_06280_),
    .X(_13579_));
 sky130_fd_sc_hd__maj3_4 _19794_ (.A(\hash.CA2.a_dash[10] ),
    .B(\hash.CA1.S0.X[10] ),
    .C(\hash.CA1.b[10] ),
    .X(_13583_));
 sky130_fd_sc_hd__o211ai_1 _19795_ (.A1(_04614_),
    .A2(_06065_),
    .B1(_06002_),
    .C1(\hash.CA2.a_dash[11] ),
    .Y(_07921_));
 sky130_fd_sc_hd__o21ai_0 _19796_ (.A1(_06066_),
    .A2(_06282_),
    .B1(_07921_),
    .Y(_13587_));
 sky130_fd_sc_hd__maj3_1 _19797_ (.A(\hash.CA2.a_dash[12] ),
    .B(\hash.CA1.S0.X[12] ),
    .C(_06283_),
    .X(_13591_));
 sky130_fd_sc_hd__a21oi_1 _19798_ (.A1(\hash.CA2.a_dash[13] ),
    .A2(_04437_),
    .B1(_06079_),
    .Y(_07922_));
 sky130_fd_sc_hd__o21ai_2 _19799_ (.A1(_04638_),
    .A2(_07922_),
    .B1(_06002_),
    .Y(_13595_));
 sky130_fd_sc_hd__a21boi_0 _19800_ (.A1(\hash.CA2.a_dash[14] ),
    .A2(_04636_),
    .B1_N(_06091_),
    .Y(_07923_));
 sky130_fd_sc_hd__o21ai_0 _19801_ (.A1(_04646_),
    .A2(_07923_),
    .B1(_06002_),
    .Y(_13599_));
 sky130_fd_sc_hd__maj3_1 _19802_ (.A(\hash.CA2.a_dash[15] ),
    .B(\hash.CA1.S0.X[15] ),
    .C(\hash.CA1.b[15] ),
    .X(_13603_));
 sky130_fd_sc_hd__maj3_4 _19803_ (.A(\hash.CA2.a_dash[16] ),
    .B(\hash.CA1.S0.X[16] ),
    .C(\hash.CA1.b[16] ),
    .X(_13607_));
 sky130_fd_sc_hd__nor2_1 _19804_ (.A(\hash.CA2.a_dash[17] ),
    .B(_04520_),
    .Y(_07924_));
 sky130_fd_sc_hd__a21oi_1 _19805_ (.A1(\hash.CA2.a_dash[17] ),
    .A2(_04520_),
    .B1(\hash.CA1.S0.X[17] ),
    .Y(_07925_));
 sky130_fd_sc_hd__o21ai_0 _19806_ (.A1(_07924_),
    .A2(_07925_),
    .B1(_06002_),
    .Y(_13611_));
 sky130_fd_sc_hd__a21oi_1 _19807_ (.A1(\hash.CA2.a_dash[18] ),
    .A2(_04541_),
    .B1(_06121_),
    .Y(_07926_));
 sky130_fd_sc_hd__o21ai_1 _19808_ (.A1(_04672_),
    .A2(_07926_),
    .B1(_06002_),
    .Y(_13615_));
 sky130_fd_sc_hd__a211oi_1 _19809_ (.A1(_04559_),
    .A2(_06132_),
    .B1(net341),
    .C1(\hash.CA2.a_dash[19] ),
    .Y(_07927_));
 sky130_fd_sc_hd__nor2_1 _19810_ (.A(\hash.CA1.S0.X[19] ),
    .B(_06284_),
    .Y(_07928_));
 sky130_fd_sc_hd__nor2_2 _19811_ (.A(_07927_),
    .B(_07928_),
    .Y(_13619_));
 sky130_fd_sc_hd__nand2_1 _19812_ (.A(_04577_),
    .B(_06148_),
    .Y(_07929_));
 sky130_fd_sc_hd__o21ai_2 _19813_ (.A1(_06148_),
    .A2(\hash.CA1.b[20] ),
    .B1(\hash.CA2.a_dash[20] ),
    .Y(_07930_));
 sky130_fd_sc_hd__nand2_4 _19814_ (.A(_07929_),
    .B(_07930_),
    .Y(_13623_));
 sky130_fd_sc_hd__a21oi_2 _19815_ (.A1(\hash.CA2.a_dash[21] ),
    .A2(_04596_),
    .B1(_06155_),
    .Y(_07931_));
 sky130_fd_sc_hd__o21ai_4 _19816_ (.A1(_04697_),
    .A2(_07931_),
    .B1(_06002_),
    .Y(_13627_));
 sky130_fd_sc_hd__nand2_1 _19817_ (.A(_04704_),
    .B(net1127),
    .Y(_07932_));
 sky130_fd_sc_hd__o21ai_2 _19818_ (.A1(\hash.CA2.a_dash[22] ),
    .A2(_04420_),
    .B1(_07932_),
    .Y(_07933_));
 sky130_fd_sc_hd__nand2_1 _19819_ (.A(_06002_),
    .B(_07933_),
    .Y(_13631_));
 sky130_fd_sc_hd__o21ai_0 _19820_ (.A1(\hash.CA1.S0.X[23] ),
    .A2(_06285_),
    .B1(\hash.CA2.a_dash[23] ),
    .Y(_07934_));
 sky130_fd_sc_hd__o21ai_2 _19821_ (.A1(_06172_),
    .A2(_06895_),
    .B1(_07934_),
    .Y(_13635_));
 sky130_fd_sc_hd__o31a_1 _19822_ (.A1(_13402_),
    .A2(_13394_),
    .A3(_06177_),
    .B1(_06178_),
    .X(_07935_));
 sky130_fd_sc_hd__o21ai_2 _19823_ (.A1(\hash.CA2.a_dash[24] ),
    .A2(_04726_),
    .B1(_07935_),
    .Y(_07936_));
 sky130_fd_sc_hd__a21oi_4 _19824_ (.A1(_04727_),
    .A2(_07936_),
    .B1(net341),
    .Y(_13639_));
 sky130_fd_sc_hd__maj3_4 _19825_ (.A(\hash.CA2.a_dash[25] ),
    .B(\hash.CA1.S0.X[25] ),
    .C(\hash.CA1.b[25] ),
    .X(_13643_));
 sky130_fd_sc_hd__maj3_2 _19826_ (.A(\hash.CA2.a_dash[26] ),
    .B(_06201_),
    .C(\hash.CA1.b[26] ),
    .X(_13647_));
 sky130_fd_sc_hd__maj3_1 _19827_ (.A(\hash.CA2.a_dash[27] ),
    .B(net1069),
    .C(_06210_),
    .X(_07937_));
 sky130_fd_sc_hd__or2_4 _19828_ (.A(net341),
    .B(_07937_),
    .X(_13651_));
 sky130_fd_sc_hd__o21ai_2 _19829_ (.A1(_06215_),
    .A2(_06217_),
    .B1(_04756_),
    .Y(_07938_));
 sky130_fd_sc_hd__o21ai_0 _19830_ (.A1(\hash.CA2.a_dash[28] ),
    .A2(_04554_),
    .B1(_07938_),
    .Y(_07939_));
 sky130_fd_sc_hd__nand2_2 _19831_ (.A(_06002_),
    .B(_07939_),
    .Y(_13655_));
 sky130_fd_sc_hd__a21oi_1 _19832_ (.A1(\hash.CA2.a_dash[29] ),
    .A2(_04754_),
    .B1(\hash.CA1.S0.X[29] ),
    .Y(_07940_));
 sky130_fd_sc_hd__o21ai_2 _19833_ (.A1(_04762_),
    .A2(_07940_),
    .B1(_06002_),
    .Y(_13659_));
 sky130_fd_sc_hd__a31oi_2 _19834_ (.A1(_04770_),
    .A2(_06232_),
    .A3(_06233_),
    .B1(_04771_),
    .Y(_07941_));
 sky130_fd_sc_hd__nor2_1 _19835_ (.A(net341),
    .B(_07941_),
    .Y(_13663_));
 sky130_fd_sc_hd__inv_1 _19836_ (.A(_12373_),
    .Y(_13667_));
 sky130_fd_sc_hd__clkinv_1 _19837_ (.A(_12369_),
    .Y(_12379_));
 sky130_fd_sc_hd__xor2_2 _19838_ (.A(_13678_),
    .B(_12380_),
    .X(\hash.CA1.p4[3] ));
 sky130_fd_sc_hd__inv_1 _19839_ (.A(_12384_),
    .Y(_13682_));
 sky130_fd_sc_hd__a21o_1 _19840_ (.A1(_12378_),
    .A2(_13672_),
    .B1(_13671_),
    .X(_07942_));
 sky130_fd_sc_hd__a21oi_2 _19841_ (.A1(_13678_),
    .A2(_07942_),
    .B1(_13677_),
    .Y(_07943_));
 sky130_fd_sc_hd__xnor2_2 _19842_ (.A(_13684_),
    .B(_07943_),
    .Y(\hash.CA1.p4[4] ));
 sky130_fd_sc_hd__a21o_1 _19843_ (.A1(_13678_),
    .A2(_12380_),
    .B1(_13677_),
    .X(_07944_));
 sky130_fd_sc_hd__a21oi_2 _19844_ (.A1(_13684_),
    .A2(_07944_),
    .B1(_13683_),
    .Y(_07945_));
 sky130_fd_sc_hd__xnor2_2 _19845_ (.A(_13690_),
    .B(_07945_),
    .Y(\hash.CA1.p4[5] ));
 sky130_fd_sc_hd__inv_1 _19846_ (.A(_12392_),
    .Y(_13694_));
 sky130_fd_sc_hd__inv_1 _19847_ (.A(_13684_),
    .Y(_07946_));
 sky130_fd_sc_hd__o21bai_1 _19848_ (.A1(_07946_),
    .A2(_07943_),
    .B1_N(_13683_),
    .Y(_07947_));
 sky130_fd_sc_hd__a21o_4 _19849_ (.A1(_13690_),
    .A2(_07947_),
    .B1(_13689_),
    .X(_07948_));
 sky130_fd_sc_hd__xor2_2 _19850_ (.A(_13696_),
    .B(_07948_),
    .X(\hash.CA1.p4[6] ));
 sky130_fd_sc_hd__inv_1 _19851_ (.A(_13690_),
    .Y(_07949_));
 sky130_fd_sc_hd__o21bai_1 _19852_ (.A1(_07949_),
    .A2(_07945_),
    .B1_N(_13689_),
    .Y(_07950_));
 sky130_fd_sc_hd__a21oi_1 _19853_ (.A1(_13696_),
    .A2(_07950_),
    .B1(_13695_),
    .Y(_07951_));
 sky130_fd_sc_hd__xnor2_1 _19854_ (.A(_13702_),
    .B(_07951_),
    .Y(\hash.CA1.p4[7] ));
 sky130_fd_sc_hd__inv_1 _19855_ (.A(_12400_),
    .Y(_13706_));
 sky130_fd_sc_hd__a21oi_2 _19856_ (.A1(_13696_),
    .A2(_07948_),
    .B1(_13695_),
    .Y(_07952_));
 sky130_fd_sc_hd__inv_1 _19857_ (.A(_07952_),
    .Y(_07953_));
 sky130_fd_sc_hd__a21oi_1 _19858_ (.A1(_13702_),
    .A2(_07953_),
    .B1(_13701_),
    .Y(_07954_));
 sky130_fd_sc_hd__xnor2_1 _19859_ (.A(_13709_),
    .B(_07954_),
    .Y(\hash.CA1.p4[8] ));
 sky130_fd_sc_hd__inv_1 _19860_ (.A(_12405_),
    .Y(_13713_));
 sky130_fd_sc_hd__nand2_2 _19861_ (.A(_13702_),
    .B(_13709_),
    .Y(_07955_));
 sky130_fd_sc_hd__a21oi_1 _19862_ (.A1(_13709_),
    .A2(_13701_),
    .B1(_13708_),
    .Y(_07956_));
 sky130_fd_sc_hd__o21ai_0 _19863_ (.A1(_07951_),
    .A2(_07955_),
    .B1(_07956_),
    .Y(_07957_));
 sky130_fd_sc_hd__xor2_1 _19864_ (.A(_13715_),
    .B(_07957_),
    .X(\hash.CA1.p4[9] ));
 sky130_fd_sc_hd__nand2b_1 _19865_ (.A_N(_13714_),
    .B(_07956_),
    .Y(_07958_));
 sky130_fd_sc_hd__o21bai_4 _19866_ (.A1(_07952_),
    .A2(_07955_),
    .B1_N(_07958_),
    .Y(_07959_));
 sky130_fd_sc_hd__o21a_4 _19867_ (.A1(_13715_),
    .A2(_13714_),
    .B1(_13720_),
    .X(_07960_));
 sky130_fd_sc_hd__o21ai_0 _19868_ (.A1(_07952_),
    .A2(_07955_),
    .B1(_07956_),
    .Y(_07961_));
 sky130_fd_sc_hd__a211oi_1 _19869_ (.A1(_13715_),
    .A2(_07961_),
    .B1(_13714_),
    .C1(_13720_),
    .Y(_07962_));
 sky130_fd_sc_hd__a21oi_2 _19870_ (.A1(_07959_),
    .A2(_07960_),
    .B1(_07962_),
    .Y(\hash.CA1.p4[10] ));
 sky130_fd_sc_hd__a211oi_1 _19871_ (.A1(_13696_),
    .A2(_07950_),
    .B1(_07958_),
    .C1(_13695_),
    .Y(_07963_));
 sky130_fd_sc_hd__a21boi_0 _19872_ (.A1(_07956_),
    .A2(_07955_),
    .B1_N(_13715_),
    .Y(_07964_));
 sky130_fd_sc_hd__o21ai_0 _19873_ (.A1(_13714_),
    .A2(_07964_),
    .B1(_13720_),
    .Y(_07965_));
 sky130_fd_sc_hd__nor2_1 _19874_ (.A(_07963_),
    .B(_07965_),
    .Y(_07966_));
 sky130_fd_sc_hd__nor2_2 _19875_ (.A(_13719_),
    .B(_07966_),
    .Y(_07967_));
 sky130_fd_sc_hd__xnor2_1 _19876_ (.A(_13726_),
    .B(_07967_),
    .Y(\hash.CA1.p4[11] ));
 sky130_fd_sc_hd__inv_2 _19877_ (.A(_12416_),
    .Y(_13730_));
 sky130_fd_sc_hd__inv_1 _19878_ (.A(_13726_),
    .Y(_07968_));
 sky130_fd_sc_hd__a21oi_1 _19879_ (.A1(_07959_),
    .A2(_07960_),
    .B1(_13719_),
    .Y(_07969_));
 sky130_fd_sc_hd__o21bai_1 _19880_ (.A1(_07968_),
    .A2(_07969_),
    .B1_N(_13725_),
    .Y(_07970_));
 sky130_fd_sc_hd__xor2_1 _19881_ (.A(_13733_),
    .B(_07970_),
    .X(\hash.CA1.p4[12] ));
 sky130_fd_sc_hd__inv_1 _19882_ (.A(_12421_),
    .Y(_13737_));
 sky130_fd_sc_hd__o21bai_1 _19883_ (.A1(_07968_),
    .A2(_07967_),
    .B1_N(_13725_),
    .Y(_07971_));
 sky130_fd_sc_hd__a21oi_1 _19884_ (.A1(_13733_),
    .A2(_07971_),
    .B1(_13732_),
    .Y(_07972_));
 sky130_fd_sc_hd__xnor2_1 _19885_ (.A(_13739_),
    .B(_07972_),
    .Y(\hash.CA1.p4[13] ));
 sky130_fd_sc_hd__a2111oi_2 _19886_ (.A1(_07959_),
    .A2(_07960_),
    .B1(_13719_),
    .C1(_13725_),
    .D1(_13732_),
    .Y(_07973_));
 sky130_fd_sc_hd__o21a_1 _19887_ (.A1(_13726_),
    .A2(_13725_),
    .B1(_13733_),
    .X(_07974_));
 sky130_fd_sc_hd__nor2_1 _19888_ (.A(_13732_),
    .B(_07974_),
    .Y(_07975_));
 sky130_fd_sc_hd__nor2_1 _19889_ (.A(_07973_),
    .B(_07975_),
    .Y(_07976_));
 sky130_fd_sc_hd__a21oi_1 _19890_ (.A1(_13739_),
    .A2(_07976_),
    .B1(_13738_),
    .Y(_07977_));
 sky130_fd_sc_hd__xnor2_1 _19891_ (.A(_13745_),
    .B(_07977_),
    .Y(\hash.CA1.p4[14] ));
 sky130_fd_sc_hd__inv_1 _19892_ (.A(_12429_),
    .Y(_13749_));
 sky130_fd_sc_hd__nand3_1 _19893_ (.A(_13726_),
    .B(_13733_),
    .C(_13739_),
    .Y(_07978_));
 sky130_fd_sc_hd__a21o_1 _19894_ (.A1(_13733_),
    .A2(_13725_),
    .B1(_13732_),
    .X(_07979_));
 sky130_fd_sc_hd__a21oi_1 _19895_ (.A1(_13739_),
    .A2(_07979_),
    .B1(_13738_),
    .Y(_07980_));
 sky130_fd_sc_hd__o21ai_0 _19896_ (.A1(_07967_),
    .A2(_07978_),
    .B1(_07980_),
    .Y(_07981_));
 sky130_fd_sc_hd__a21oi_1 _19897_ (.A1(_13745_),
    .A2(_07981_),
    .B1(_13744_),
    .Y(_07982_));
 sky130_fd_sc_hd__xnor2_1 _19898_ (.A(_13752_),
    .B(_07982_),
    .Y(\hash.CA1.p4[15] ));
 sky130_fd_sc_hd__inv_1 _19899_ (.A(_12434_),
    .Y(_13756_));
 sky130_fd_sc_hd__and2_4 _19900_ (.A(_13745_),
    .B(_13752_),
    .X(_07983_));
 sky130_fd_sc_hd__o211ai_1 _19901_ (.A1(_13732_),
    .A2(_07974_),
    .B1(_07983_),
    .C1(_13739_),
    .Y(_07984_));
 sky130_fd_sc_hd__a22oi_1 _19902_ (.A1(_13752_),
    .A2(_13744_),
    .B1(_07983_),
    .B2(_13738_),
    .Y(_07985_));
 sky130_fd_sc_hd__nor2b_1 _19903_ (.A(_13751_),
    .B_N(_07985_),
    .Y(_07986_));
 sky130_fd_sc_hd__o21ai_0 _19904_ (.A1(_07973_),
    .A2(_07984_),
    .B1(_07986_),
    .Y(_07987_));
 sky130_fd_sc_hd__xor2_1 _19905_ (.A(_13759_),
    .B(_07987_),
    .X(\hash.CA1.p4[16] ));
 sky130_fd_sc_hd__inv_1 _19906_ (.A(_12439_),
    .Y(_13763_));
 sky130_fd_sc_hd__nor3_1 _19907_ (.A(_07963_),
    .B(_07965_),
    .C(_07978_),
    .Y(_07988_));
 sky130_fd_sc_hd__inv_1 _19908_ (.A(_13719_),
    .Y(_07989_));
 sky130_fd_sc_hd__o21ai_0 _19909_ (.A1(_07989_),
    .A2(_07978_),
    .B1(_07980_),
    .Y(_07990_));
 sky130_fd_sc_hd__o211ai_1 _19910_ (.A1(_07988_),
    .A2(_07990_),
    .B1(_07983_),
    .C1(_13759_),
    .Y(_07991_));
 sky130_fd_sc_hd__and3_1 _19911_ (.A(_13752_),
    .B(_13759_),
    .C(_13744_),
    .X(_07992_));
 sky130_fd_sc_hd__a21oi_1 _19912_ (.A1(_13759_),
    .A2(_13751_),
    .B1(_07992_),
    .Y(_07993_));
 sky130_fd_sc_hd__nand3b_1 _19913_ (.A_N(_13758_),
    .B(_07991_),
    .C(_07993_),
    .Y(_07994_));
 sky130_fd_sc_hd__xor2_1 _19914_ (.A(_13766_),
    .B(_07994_),
    .X(\hash.CA1.p4[17] ));
 sky130_fd_sc_hd__inv_1 _19915_ (.A(_12444_),
    .Y(_13770_));
 sky130_fd_sc_hd__nor3_1 _19916_ (.A(_13751_),
    .B(_13758_),
    .C(_13765_),
    .Y(_07995_));
 sky130_fd_sc_hd__o211ai_1 _19917_ (.A1(_07973_),
    .A2(_07984_),
    .B1(_07985_),
    .C1(_07995_),
    .Y(_07996_));
 sky130_fd_sc_hd__or2_0 _19918_ (.A(_13766_),
    .B(_13765_),
    .X(_07997_));
 sky130_fd_sc_hd__o31a_1 _19919_ (.A1(_13759_),
    .A2(_13758_),
    .A3(_13765_),
    .B1(_07997_),
    .X(_07998_));
 sky130_fd_sc_hd__nand2_2 _19920_ (.A(_07996_),
    .B(_07998_),
    .Y(_07999_));
 sky130_fd_sc_hd__xnor2_1 _19921_ (.A(_13772_),
    .B(_07999_),
    .Y(\hash.CA1.p4[18] ));
 sky130_fd_sc_hd__nor3_1 _19922_ (.A(_13758_),
    .B(_13765_),
    .C(_13771_),
    .Y(_08000_));
 sky130_fd_sc_hd__a21oi_1 _19923_ (.A1(_13772_),
    .A2(_07997_),
    .B1(_13771_),
    .Y(_08001_));
 sky130_fd_sc_hd__a31oi_2 _19924_ (.A1(_07991_),
    .A2(_07993_),
    .A3(_08000_),
    .B1(_08001_),
    .Y(_08002_));
 sky130_fd_sc_hd__xor2_1 _19925_ (.A(_13777_),
    .B(_08002_),
    .X(\hash.CA1.p4[19] ));
 sky130_fd_sc_hd__nand3_1 _19926_ (.A(_13772_),
    .B(_13777_),
    .C(_13782_),
    .Y(_08003_));
 sky130_fd_sc_hd__and3_1 _19927_ (.A(_13777_),
    .B(_13782_),
    .C(_13771_),
    .X(_08004_));
 sky130_fd_sc_hd__a21oi_1 _19928_ (.A1(_13782_),
    .A2(_13776_),
    .B1(_08004_),
    .Y(_08005_));
 sky130_fd_sc_hd__o21ai_2 _19929_ (.A1(_07999_),
    .A2(_08003_),
    .B1(_08005_),
    .Y(_08006_));
 sky130_fd_sc_hd__a31o_1 _19930_ (.A1(_13772_),
    .A2(_07996_),
    .A3(_07998_),
    .B1(_13771_),
    .X(_08007_));
 sky130_fd_sc_hd__a211oi_1 _19931_ (.A1(_13777_),
    .A2(_08007_),
    .B1(_13776_),
    .C1(_13782_),
    .Y(_08008_));
 sky130_fd_sc_hd__nor2_1 _19932_ (.A(_08006_),
    .B(_08008_),
    .Y(\hash.CA1.p4[20] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_984 ();
 sky130_fd_sc_hd__a21o_1 _19934_ (.A1(_13777_),
    .A2(_08002_),
    .B1(_13776_),
    .X(_08010_));
 sky130_fd_sc_hd__a21oi_1 _19935_ (.A1(_13782_),
    .A2(_08010_),
    .B1(_13781_),
    .Y(_08011_));
 sky130_fd_sc_hd__xnor2_1 _19936_ (.A(_13787_),
    .B(_08011_),
    .Y(\hash.CA1.p4[21] ));
 sky130_fd_sc_hd__inv_1 _19937_ (.A(_13781_),
    .Y(_08012_));
 sky130_fd_sc_hd__o211ai_1 _19938_ (.A1(_07999_),
    .A2(_08003_),
    .B1(_08005_),
    .C1(_08012_),
    .Y(_08013_));
 sky130_fd_sc_hd__a21oi_1 _19939_ (.A1(_13787_),
    .A2(_08013_),
    .B1(_13786_),
    .Y(_08014_));
 sky130_fd_sc_hd__xnor2_1 _19940_ (.A(_13792_),
    .B(_08014_),
    .Y(\hash.CA1.p4[22] ));
 sky130_fd_sc_hd__and3_1 _19941_ (.A(_13777_),
    .B(_13782_),
    .C(_13787_),
    .X(_08015_));
 sky130_fd_sc_hd__nand2_1 _19942_ (.A(_13787_),
    .B(_13781_),
    .Y(_08016_));
 sky130_fd_sc_hd__nand3_1 _19943_ (.A(_13782_),
    .B(_13787_),
    .C(_13776_),
    .Y(_08017_));
 sky130_fd_sc_hd__nand2_1 _19944_ (.A(_08016_),
    .B(_08017_),
    .Y(_08018_));
 sky130_fd_sc_hd__a211o_1 _19945_ (.A1(_08002_),
    .A2(_08015_),
    .B1(_08018_),
    .C1(_13786_),
    .X(_08019_));
 sky130_fd_sc_hd__a21o_4 _19946_ (.A1(_13792_),
    .A2(_08019_),
    .B1(_13791_),
    .X(_08020_));
 sky130_fd_sc_hd__xor2_1 _19947_ (.A(_13798_),
    .B(_08020_),
    .X(\hash.CA1.p4[23] ));
 sky130_fd_sc_hd__inv_1 _19948_ (.A(_12464_),
    .Y(_13802_));
 sky130_fd_sc_hd__a21o_4 _19949_ (.A1(_13798_),
    .A2(_13791_),
    .B1(_13797_),
    .X(_08021_));
 sky130_fd_sc_hd__nand2_1 _19950_ (.A(_13792_),
    .B(_13798_),
    .Y(_08022_));
 sky130_fd_sc_hd__nor2_1 _19951_ (.A(_13787_),
    .B(_13786_),
    .Y(_08023_));
 sky130_fd_sc_hd__o21bai_1 _19952_ (.A1(_08022_),
    .A2(_08023_),
    .B1_N(_08021_),
    .Y(_08024_));
 sky130_fd_sc_hd__o41ai_2 _19953_ (.A1(_13781_),
    .A2(_13786_),
    .A3(_08006_),
    .A4(_08021_),
    .B1(_08024_),
    .Y(_08025_));
 sky130_fd_sc_hd__xnor2_1 _19954_ (.A(_13805_),
    .B(_08025_),
    .Y(\hash.CA1.p4[24] ));
 sky130_fd_sc_hd__inv_1 _19955_ (.A(_12469_),
    .Y(_13809_));
 sky130_fd_sc_hd__clkinv_1 _19956_ (.A(_13812_),
    .Y(_08026_));
 sky130_fd_sc_hd__a21oi_1 _19957_ (.A1(_13805_),
    .A2(_13797_),
    .B1(_13804_),
    .Y(_08027_));
 sky130_fd_sc_hd__nand3_1 _19958_ (.A(_13798_),
    .B(_13805_),
    .C(_08020_),
    .Y(_08028_));
 sky130_fd_sc_hd__nand2_1 _19959_ (.A(_08027_),
    .B(_08028_),
    .Y(_08029_));
 sky130_fd_sc_hd__xnor2_1 _19960_ (.A(_08026_),
    .B(_08029_),
    .Y(\hash.CA1.p4[25] ));
 sky130_fd_sc_hd__inv_1 _19961_ (.A(_12474_),
    .Y(_13816_));
 sky130_fd_sc_hd__nor2_1 _19962_ (.A(_08014_),
    .B(_08022_),
    .Y(_08030_));
 sky130_fd_sc_hd__a21oi_1 _19963_ (.A1(_13805_),
    .A2(_08021_),
    .B1(_13804_),
    .Y(_08031_));
 sky130_fd_sc_hd__o21bai_1 _19964_ (.A1(_08026_),
    .A2(_08031_),
    .B1_N(_13811_),
    .Y(_08032_));
 sky130_fd_sc_hd__a31oi_1 _19965_ (.A1(_13805_),
    .A2(_13812_),
    .A3(_08030_),
    .B1(_08032_),
    .Y(_08033_));
 sky130_fd_sc_hd__xnor2_2 _19966_ (.A(_13819_),
    .B(_08033_),
    .Y(\hash.CA1.p4[26] ));
 sky130_fd_sc_hd__inv_1 _19967_ (.A(_12479_),
    .Y(_13823_));
 sky130_fd_sc_hd__inv_2 _19968_ (.A(_13826_),
    .Y(_08034_));
 sky130_fd_sc_hd__nand2_2 _19969_ (.A(_13798_),
    .B(_08020_),
    .Y(_08035_));
 sky130_fd_sc_hd__nand3_2 _19970_ (.A(_13805_),
    .B(_13812_),
    .C(_13819_),
    .Y(_08036_));
 sky130_fd_sc_hd__o21bai_1 _19971_ (.A1(_08026_),
    .A2(_08027_),
    .B1_N(_13811_),
    .Y(_08037_));
 sky130_fd_sc_hd__a21oi_1 _19972_ (.A1(_13819_),
    .A2(_08037_),
    .B1(_13818_),
    .Y(_08038_));
 sky130_fd_sc_hd__o21ai_2 _19973_ (.A1(_08035_),
    .A2(_08036_),
    .B1(_08038_),
    .Y(_08039_));
 sky130_fd_sc_hd__xnor2_1 _19974_ (.A(_08034_),
    .B(_08039_),
    .Y(\hash.CA1.p4[27] ));
 sky130_fd_sc_hd__inv_1 _19975_ (.A(_12484_),
    .Y(_13830_));
 sky130_fd_sc_hd__a21o_1 _19976_ (.A1(_13812_),
    .A2(_13804_),
    .B1(_13811_),
    .X(_08040_));
 sky130_fd_sc_hd__a21oi_1 _19977_ (.A1(_13819_),
    .A2(_08040_),
    .B1(_13818_),
    .Y(_08041_));
 sky130_fd_sc_hd__o21ai_0 _19978_ (.A1(_08025_),
    .A2(_08036_),
    .B1(_08041_),
    .Y(_08042_));
 sky130_fd_sc_hd__a21oi_1 _19979_ (.A1(_13826_),
    .A2(_08042_),
    .B1(_13825_),
    .Y(_08043_));
 sky130_fd_sc_hd__xnor2_1 _19980_ (.A(_13833_),
    .B(_08043_),
    .Y(\hash.CA1.p4[28] ));
 sky130_fd_sc_hd__clkinv_1 _19981_ (.A(_12489_),
    .Y(_13837_));
 sky130_fd_sc_hd__a21o_1 _19982_ (.A1(_13826_),
    .A2(_08039_),
    .B1(_13825_),
    .X(_08044_));
 sky130_fd_sc_hd__a21oi_1 _19983_ (.A1(_13833_),
    .A2(_08044_),
    .B1(_13832_),
    .Y(_08045_));
 sky130_fd_sc_hd__xnor2_1 _19984_ (.A(_13839_),
    .B(_08045_),
    .Y(\hash.CA1.p4[29] ));
 sky130_fd_sc_hd__a21oi_1 _19985_ (.A1(_13819_),
    .A2(_08032_),
    .B1(_13818_),
    .Y(_08046_));
 sky130_fd_sc_hd__nor2_1 _19986_ (.A(_08034_),
    .B(_08046_),
    .Y(_08047_));
 sky130_fd_sc_hd__o21a_1 _19987_ (.A1(_13825_),
    .A2(_08047_),
    .B1(_13833_),
    .X(_08048_));
 sky130_fd_sc_hd__o21ai_1 _19988_ (.A1(_13832_),
    .A2(_08048_),
    .B1(_13839_),
    .Y(_08049_));
 sky130_fd_sc_hd__nand2_1 _19989_ (.A(_13833_),
    .B(_13839_),
    .Y(_08050_));
 sky130_fd_sc_hd__or3_4 _19990_ (.A(_08034_),
    .B(_08036_),
    .C(_08050_),
    .X(_08051_));
 sky130_fd_sc_hd__nor2_1 _19991_ (.A(_08022_),
    .B(_08051_),
    .Y(_08052_));
 sky130_fd_sc_hd__nand2b_1 _19992_ (.A_N(_13786_),
    .B(_08016_),
    .Y(_08053_));
 sky130_fd_sc_hd__a21oi_1 _19993_ (.A1(_08052_),
    .A2(_08053_),
    .B1(_13838_),
    .Y(_08054_));
 sky130_fd_sc_hd__nand3_1 _19994_ (.A(_13787_),
    .B(_08006_),
    .C(_08052_),
    .Y(_08055_));
 sky130_fd_sc_hd__nand3_2 _19995_ (.A(_08049_),
    .B(_08054_),
    .C(_08055_),
    .Y(_08056_));
 sky130_fd_sc_hd__xor2_1 _19996_ (.A(_13844_),
    .B(_08056_),
    .X(\hash.CA1.p4[30] ));
 sky130_fd_sc_hd__xnor2_1 _19997_ (.A(\hash.CA1.S1.X[6] ),
    .B(_06575_),
    .Y(_08057_));
 sky130_fd_sc_hd__xnor2_2 _19998_ (.A(_06683_),
    .B(_08057_),
    .Y(_13861_));
 sky130_fd_sc_hd__xor2_1 _19999_ (.A(\hash.CA1.S1.X[7] ),
    .B(_06581_),
    .X(_08058_));
 sky130_fd_sc_hd__xnor2_1 _20000_ (.A(_06689_),
    .B(_08058_),
    .Y(_12501_));
 sky130_fd_sc_hd__xnor2_1 _20001_ (.A(_06552_),
    .B(\hash.CA1.S1.X[13] ),
    .Y(_08059_));
 sky130_fd_sc_hd__xnor2_1 _20002_ (.A(_06699_),
    .B(_08059_),
    .Y(_13869_));
 sky130_fd_sc_hd__xnor2_1 _20003_ (.A(_06559_),
    .B(_06597_),
    .Y(_08060_));
 sky130_fd_sc_hd__xnor2_2 _20004_ (.A(_06707_),
    .B(_08060_),
    .Y(_13877_));
 sky130_fd_sc_hd__xnor2_1 _20005_ (.A(\hash.CA1.S1.X[10] ),
    .B(_06610_),
    .Y(_08061_));
 sky130_fd_sc_hd__xnor2_4 _20006_ (.A(\hash.CA1.S1.X[29] ),
    .B(_08061_),
    .Y(_13886_));
 sky130_fd_sc_hd__inv_1 _20007_ (.A(_12516_),
    .Y(_13890_));
 sky130_fd_sc_hd__nand3b_1 _20008_ (.A_N(_13884_),
    .B(_06942_),
    .C(_06943_),
    .Y(_08062_));
 sky130_fd_sc_hd__xor2_2 _20009_ (.A(_13895_),
    .B(_08062_),
    .X(_12524_));
 sky130_fd_sc_hd__xnor2_1 _20010_ (.A(_06575_),
    .B(\hash.CA1.S1.X[16] ),
    .Y(_08063_));
 sky130_fd_sc_hd__xnor2_2 _20011_ (.A(_08063_),
    .B(\hash.CA1.S1.X[30] ),
    .Y(_13896_));
 sky130_fd_sc_hd__inv_1 _20012_ (.A(_12521_),
    .Y(_13900_));
 sky130_fd_sc_hd__xnor2_1 _20013_ (.A(_06581_),
    .B(_06624_),
    .Y(_08064_));
 sky130_fd_sc_hd__xnor2_1 _20014_ (.A(\hash.CA1.S1.X[31] ),
    .B(_08064_),
    .Y(_13905_));
 sky130_fd_sc_hd__nor2_1 _20015_ (.A(\hash.CA1.S1.X[0] ),
    .B(\hash.CA1.S1.X[13] ),
    .Y(_08065_));
 sky130_fd_sc_hd__a21oi_2 _20016_ (.A1(_13445_),
    .A2(\hash.CA1.S1.X[13] ),
    .B1(_08065_),
    .Y(_08066_));
 sky130_fd_sc_hd__xnor2_1 _20017_ (.A(_06634_),
    .B(_08066_),
    .Y(_13913_));
 sky130_fd_sc_hd__nor2_1 _20018_ (.A(\hash.CA1.S1.X[1] ),
    .B(_06642_),
    .Y(_08067_));
 sky130_fd_sc_hd__a21oi_1 _20019_ (.A1(_12365_),
    .A2(_06642_),
    .B1(_08067_),
    .Y(_08068_));
 sky130_fd_sc_hd__xnor2_2 _20020_ (.A(\hash.CA1.S1.X[14] ),
    .B(_08068_),
    .Y(_13921_));
 sky130_fd_sc_hd__xnor2_1 _20021_ (.A(\hash.CA1.S1.X[2] ),
    .B(_06610_),
    .Y(_08069_));
 sky130_fd_sc_hd__xnor2_1 _20022_ (.A(\hash.CA1.S1.X[20] ),
    .B(_08069_),
    .Y(_13930_));
 sky130_fd_sc_hd__xnor2_2 _20023_ (.A(_07117_),
    .B(_13933_),
    .Y(_12543_));
 sky130_fd_sc_hd__clkinv_1 _20024_ (.A(_12541_),
    .Y(_13934_));
 sky130_fd_sc_hd__xnor2_1 _20025_ (.A(\hash.CA1.S1.X[3] ),
    .B(\hash.CA1.S1.X[16] ),
    .Y(_08070_));
 sky130_fd_sc_hd__xnor2_1 _20026_ (.A(\hash.CA1.S1.X[21] ),
    .B(_08070_),
    .Y(_13939_));
 sky130_fd_sc_hd__xnor2_1 _20027_ (.A(_06524_),
    .B(_06624_),
    .Y(_08071_));
 sky130_fd_sc_hd__xnor2_1 _20028_ (.A(\hash.CA1.S1.X[22] ),
    .B(_08071_),
    .Y(_13948_));
 sky130_fd_sc_hd__clkinv_1 _20029_ (.A(_12551_),
    .Y(_13952_));
 sky130_fd_sc_hd__a21oi_1 _20030_ (.A1(_06956_),
    .A2(_06971_),
    .B1(_06974_),
    .Y(_08072_));
 sky130_fd_sc_hd__o21ai_1 _20031_ (.A1(_06969_),
    .A2(_08072_),
    .B1(_07002_),
    .Y(_08073_));
 sky130_fd_sc_hd__xnor2_2 _20032_ (.A(_06982_),
    .B(_08073_),
    .Y(_12559_));
 sky130_fd_sc_hd__xnor2_1 _20033_ (.A(_06531_),
    .B(_06634_),
    .Y(_08074_));
 sky130_fd_sc_hd__xnor2_1 _20034_ (.A(\hash.CA1.S1.X[23] ),
    .B(_08074_),
    .Y(_13958_));
 sky130_fd_sc_hd__xnor2_2 _20035_ (.A(_13961_),
    .B(_07119_),
    .Y(_12558_));
 sky130_fd_sc_hd__clkinv_1 _20036_ (.A(_12556_),
    .Y(_13962_));
 sky130_fd_sc_hd__a21oi_1 _20037_ (.A1(_07001_),
    .A2(_07003_),
    .B1(_13956_),
    .Y(_08075_));
 sky130_fd_sc_hd__xnor2_2 _20038_ (.A(_13966_),
    .B(_08075_),
    .Y(_12564_));
 sky130_fd_sc_hd__xnor2_1 _20039_ (.A(\hash.CA1.S1.X[6] ),
    .B(_06642_),
    .Y(_08076_));
 sky130_fd_sc_hd__xnor2_1 _20040_ (.A(_06673_),
    .B(_08076_),
    .Y(_13967_));
 sky130_fd_sc_hd__o31a_1 _20041_ (.A1(_13970_),
    .A2(_06989_),
    .A3(_07120_),
    .B1(_07012_),
    .X(_12563_));
 sky130_fd_sc_hd__xnor2_1 _20042_ (.A(\hash.CA1.S1.X[7] ),
    .B(\hash.CA1.S1.X[20] ),
    .Y(_08077_));
 sky130_fd_sc_hd__xnor2_1 _20043_ (.A(_06683_),
    .B(_08077_),
    .Y(_13975_));
 sky130_fd_sc_hd__xnor2_1 _20044_ (.A(_06552_),
    .B(\hash.CA1.S1.X[21] ),
    .Y(_08078_));
 sky130_fd_sc_hd__xnor2_1 _20045_ (.A(_06689_),
    .B(_08078_),
    .Y(_13984_));
 sky130_fd_sc_hd__clkinv_1 _20046_ (.A(_12571_),
    .Y(_13988_));
 sky130_fd_sc_hd__a21oi_1 _20047_ (.A1(_13983_),
    .A2(_07024_),
    .B1(_13982_),
    .Y(_08079_));
 sky130_fd_sc_hd__xnor2_1 _20048_ (.A(_13993_),
    .B(_08079_),
    .Y(_12579_));
 sky130_fd_sc_hd__xnor2_1 _20049_ (.A(\hash.CA1.S1.X[9] ),
    .B(\hash.CA1.S1.X[22] ),
    .Y(_08080_));
 sky130_fd_sc_hd__xnor2_1 _20050_ (.A(net1124),
    .B(_08080_),
    .Y(_13994_));
 sky130_fd_sc_hd__xnor2_1 _20051_ (.A(_13997_),
    .B(_07055_),
    .Y(_12578_));
 sky130_fd_sc_hd__clkinv_1 _20052_ (.A(_12576_),
    .Y(_13998_));
 sky130_fd_sc_hd__a31oi_1 _20053_ (.A1(_13983_),
    .A2(_13993_),
    .A3(_07008_),
    .B1(_07019_),
    .Y(_08081_));
 sky130_fd_sc_hd__xnor2_1 _20054_ (.A(_14002_),
    .B(_08081_),
    .Y(_12584_));
 sky130_fd_sc_hd__xnor2_1 _20055_ (.A(\hash.CA1.S1.X[10] ),
    .B(\hash.CA1.S1.X[23] ),
    .Y(_08082_));
 sky130_fd_sc_hd__xnor2_1 _20056_ (.A(_06707_),
    .B(_08082_),
    .Y(_14003_));
 sky130_fd_sc_hd__a21oi_1 _20057_ (.A1(_07121_),
    .A2(_07122_),
    .B1(_07041_),
    .Y(_12583_));
 sky130_fd_sc_hd__a31o_1 _20058_ (.A1(_13983_),
    .A2(_13993_),
    .A3(_07024_),
    .B1(_07019_),
    .X(_08083_));
 sky130_fd_sc_hd__a21oi_1 _20059_ (.A1(_14002_),
    .A2(_08083_),
    .B1(_14001_),
    .Y(_08084_));
 sky130_fd_sc_hd__xnor2_2 _20060_ (.A(_14010_),
    .B(_08084_),
    .Y(_12589_));
 sky130_fd_sc_hd__xnor3_1 _20061_ (.A(_06575_),
    .B(_06673_),
    .C(\hash.CA1.S1.X[29] ),
    .X(_14011_));
 sky130_fd_sc_hd__xnor2_1 _20062_ (.A(_14014_),
    .B(_07123_),
    .Y(_12588_));
 sky130_fd_sc_hd__xnor2_1 _20063_ (.A(_14018_),
    .B(_07030_),
    .Y(_12594_));
 sky130_fd_sc_hd__xnor2_1 _20064_ (.A(\hash.CA1.S1.X[12] ),
    .B(_06683_),
    .Y(_08085_));
 sky130_fd_sc_hd__xnor2_1 _20065_ (.A(net1040),
    .B(_08085_),
    .Y(_14019_));
 sky130_fd_sc_hd__xnor2_1 _20066_ (.A(_14022_),
    .B(_07125_),
    .Y(_12593_));
 sky130_fd_sc_hd__xnor2_1 _20067_ (.A(\hash.CA1.S1.X[13] ),
    .B(_06689_),
    .Y(_08086_));
 sky130_fd_sc_hd__xnor2_1 _20068_ (.A(\hash.CA1.S1.X[31] ),
    .B(_08086_),
    .Y(_14027_));
 sky130_fd_sc_hd__xnor2_1 _20069_ (.A(_14030_),
    .B(_07128_),
    .Y(_12598_));
 sky130_fd_sc_hd__nor2_1 _20070_ (.A(\hash.CA1.S1.X[0] ),
    .B(_06699_),
    .Y(_08087_));
 sky130_fd_sc_hd__a21oi_1 _20071_ (.A1(_13445_),
    .A2(_06699_),
    .B1(_08087_),
    .Y(_08088_));
 sky130_fd_sc_hd__xnor2_1 _20072_ (.A(_06597_),
    .B(_08088_),
    .Y(_14035_));
 sky130_fd_sc_hd__mux2i_1 _20073_ (.A0(_12365_),
    .A1(_13854_),
    .S(_06707_),
    .Y(_08089_));
 sky130_fd_sc_hd__xnor2_1 _20074_ (.A(_06610_),
    .B(_08089_),
    .Y(_14044_));
 sky130_fd_sc_hd__inv_1 _20075_ (.A(_12606_),
    .Y(_14048_));
 sky130_fd_sc_hd__xnor2_1 _20076_ (.A(_06514_),
    .B(\hash.CA1.S1.X[16] ),
    .Y(_08090_));
 sky130_fd_sc_hd__xnor2_1 _20077_ (.A(_06712_),
    .B(_08090_),
    .Y(_14054_));
 sky130_fd_sc_hd__inv_2 _20078_ (.A(_12611_),
    .Y(_14058_));
 sky130_fd_sc_hd__xor2_1 _20079_ (.A(\hash.CA1.S1.X[3] ),
    .B(_06624_),
    .X(_08091_));
 sky130_fd_sc_hd__xnor2_1 _20080_ (.A(net1041),
    .B(_08091_),
    .Y(_14064_));
 sky130_fd_sc_hd__inv_2 _20081_ (.A(_12616_),
    .Y(_14068_));
 sky130_fd_sc_hd__xnor2_1 _20082_ (.A(_06524_),
    .B(_06634_),
    .Y(_08092_));
 sky130_fd_sc_hd__xnor2_2 _20083_ (.A(\hash.CA1.S1.X[31] ),
    .B(_08092_),
    .Y(_14074_));
 sky130_fd_sc_hd__inv_2 _20084_ (.A(_12621_),
    .Y(_14078_));
 sky130_fd_sc_hd__nor2_1 _20085_ (.A(_14072_),
    .B(_07093_),
    .Y(_08093_));
 sky130_fd_sc_hd__xnor2_2 _20086_ (.A(_14083_),
    .B(_08093_),
    .Y(_12629_));
 sky130_fd_sc_hd__nand2_8 _20087_ (.A(_06528_),
    .B(_06530_),
    .Y(_08094_));
 sky130_fd_sc_hd__xnor2_1 _20088_ (.A(_13445_),
    .B(_08094_),
    .Y(_08095_));
 sky130_fd_sc_hd__and2_0 _20089_ (.A(_06002_),
    .B(_08095_),
    .X(_08096_));
 sky130_fd_sc_hd__xnor2_1 _20090_ (.A(_06642_),
    .B(_08096_),
    .Y(_14084_));
 sky130_fd_sc_hd__xor2_1 _20091_ (.A(_14087_),
    .B(_07129_),
    .X(_12628_));
 sky130_fd_sc_hd__inv_1 _20092_ (.A(_12626_),
    .Y(_14088_));
 sky130_fd_sc_hd__mux2i_1 _20093_ (.A0(_12365_),
    .A1(_13854_),
    .S(\hash.CA1.S1.X[6] ),
    .Y(_08097_));
 sky130_fd_sc_hd__xnor2_1 _20094_ (.A(\hash.CA1.S1.X[20] ),
    .B(_08097_),
    .Y(_14093_));
 sky130_fd_sc_hd__xnor2_1 _20095_ (.A(\hash.CA1.S1.X[2] ),
    .B(\hash.CA1.S1.X[7] ),
    .Y(_08098_));
 sky130_fd_sc_hd__xnor2_2 _20096_ (.A(\hash.CA1.S1.X[21] ),
    .B(_08098_),
    .Y(_14102_));
 sky130_fd_sc_hd__inv_1 _20097_ (.A(_12636_),
    .Y(_14106_));
 sky130_fd_sc_hd__nor3_1 _20098_ (.A(_14072_),
    .B(_14082_),
    .C(_14091_),
    .Y(_08099_));
 sky130_fd_sc_hd__nand2_1 _20099_ (.A(_14101_),
    .B(_07095_),
    .Y(_08100_));
 sky130_fd_sc_hd__a21oi_1 _20100_ (.A1(_07084_),
    .A2(_08099_),
    .B1(_08100_),
    .Y(_08101_));
 sky130_fd_sc_hd__nor2_1 _20101_ (.A(_14100_),
    .B(_08101_),
    .Y(_08102_));
 sky130_fd_sc_hd__xnor2_2 _20102_ (.A(_14111_),
    .B(_08102_),
    .Y(_12644_));
 sky130_fd_sc_hd__xnor2_1 _20103_ (.A(\hash.CA1.S1.X[3] ),
    .B(_06552_),
    .Y(_08103_));
 sky130_fd_sc_hd__xnor2_1 _20104_ (.A(\hash.CA1.S1.X[22] ),
    .B(_08103_),
    .Y(_14112_));
 sky130_fd_sc_hd__xnor2_1 _20105_ (.A(_14115_),
    .B(_07134_),
    .Y(_12643_));
 sky130_fd_sc_hd__inv_1 _20106_ (.A(_12641_),
    .Y(_14116_));
 sky130_fd_sc_hd__or3_4 _20107_ (.A(_07107_),
    .B(_07109_),
    .C(_07110_),
    .X(_12870_));
 sky130_fd_sc_hd__xnor2_1 _20108_ (.A(_06524_),
    .B(_06559_),
    .Y(_08104_));
 sky130_fd_sc_hd__xnor2_1 _20109_ (.A(\hash.CA1.S1.X[23] ),
    .B(_08104_),
    .Y(_14121_));
 sky130_fd_sc_hd__inv_1 _20110_ (.A(_12663_),
    .Y(_14128_));
 sky130_fd_sc_hd__inv_1 _20111_ (.A(_12672_),
    .Y(_14132_));
 sky130_fd_sc_hd__clkinv_1 _20112_ (.A(_12677_),
    .Y(_14136_));
 sky130_fd_sc_hd__clkinv_1 _20113_ (.A(_12682_),
    .Y(_14140_));
 sky130_fd_sc_hd__clkinv_1 _20114_ (.A(_12689_),
    .Y(_14144_));
 sky130_fd_sc_hd__clkinv_1 _20115_ (.A(_12698_),
    .Y(_14148_));
 sky130_fd_sc_hd__inv_1 _20116_ (.A(_12706_),
    .Y(_14152_));
 sky130_fd_sc_hd__clkinv_1 _20117_ (.A(_12709_),
    .Y(_12718_));
 sky130_fd_sc_hd__inv_1 _20118_ (.A(_12711_),
    .Y(_14156_));
 sky130_fd_sc_hd__inv_1 _20119_ (.A(_12716_),
    .Y(_12726_));
 sky130_fd_sc_hd__inv_1 _20120_ (.A(_12753_),
    .Y(_12762_));
 sky130_fd_sc_hd__inv_1 _20121_ (.A(_12760_),
    .Y(_12770_));
 sky130_fd_sc_hd__inv_1 _20122_ (.A(_12795_),
    .Y(_12806_));
 sky130_fd_sc_hd__inv_1 _20123_ (.A(_12811_),
    .Y(_12822_));
 sky130_fd_sc_hd__inv_1 _20124_ (.A(_12827_),
    .Y(_12838_));
 sky130_fd_sc_hd__clkinv_1 _20125_ (.A(_06782_),
    .Y(_12842_));
 sky130_fd_sc_hd__a21oi_1 _20126_ (.A1(\hash.CA2.a_dash[0] ),
    .A2(_13235_),
    .B1(_12922_),
    .Y(_08105_));
 sky130_fd_sc_hd__nor2_1 _20127_ (.A(\hash.CA2.a_dash[0] ),
    .B(_13235_),
    .Y(_08106_));
 sky130_fd_sc_hd__o21ai_0 _20128_ (.A1(_08105_),
    .A2(_08106_),
    .B1(_06002_),
    .Y(_14202_));
 sky130_fd_sc_hd__clkinvlp_4 _20129_ (.A(\count_hash2[2] ),
    .Y(_12900_));
 sky130_fd_sc_hd__clkinvlp_4 _20130_ (.A(\count_hash1[2] ),
    .Y(_12910_));
 sky130_fd_sc_hd__inv_1 _20131_ (.A(_11583_),
    .Y(_12984_));
 sky130_fd_sc_hd__inv_1 _20132_ (.A(_11591_),
    .Y(_12987_));
 sky130_fd_sc_hd__inv_1 _20133_ (.A(_11599_),
    .Y(_12991_));
 sky130_fd_sc_hd__inv_1 _20134_ (.A(_11610_),
    .Y(_12995_));
 sky130_fd_sc_hd__inv_1 _20135_ (.A(_11618_),
    .Y(_12999_));
 sky130_fd_sc_hd__inv_1 _20136_ (.A(_11626_),
    .Y(_13003_));
 sky130_fd_sc_hd__inv_1 _20137_ (.A(_11634_),
    .Y(_13007_));
 sky130_fd_sc_hd__inv_1 _20138_ (.A(_11642_),
    .Y(_13011_));
 sky130_fd_sc_hd__inv_1 _20139_ (.A(_11650_),
    .Y(_13015_));
 sky130_fd_sc_hd__inv_1 _20140_ (.A(_11658_),
    .Y(_13019_));
 sky130_fd_sc_hd__inv_1 _20141_ (.A(_11666_),
    .Y(_13023_));
 sky130_fd_sc_hd__inv_1 _20142_ (.A(_11674_),
    .Y(_13027_));
 sky130_fd_sc_hd__inv_1 _20143_ (.A(_11682_),
    .Y(_13031_));
 sky130_fd_sc_hd__inv_1 _20144_ (.A(_11690_),
    .Y(_13035_));
 sky130_fd_sc_hd__inv_1 _20145_ (.A(_11698_),
    .Y(_13039_));
 sky130_fd_sc_hd__inv_1 _20146_ (.A(_11706_),
    .Y(_13043_));
 sky130_fd_sc_hd__inv_1 _20147_ (.A(_11714_),
    .Y(_13047_));
 sky130_fd_sc_hd__inv_1 _20148_ (.A(_11722_),
    .Y(_13051_));
 sky130_fd_sc_hd__inv_1 _20149_ (.A(_11730_),
    .Y(_13055_));
 sky130_fd_sc_hd__inv_1 _20150_ (.A(_11738_),
    .Y(_13059_));
 sky130_fd_sc_hd__inv_1 _20151_ (.A(_11746_),
    .Y(_13063_));
 sky130_fd_sc_hd__inv_1 _20152_ (.A(_11754_),
    .Y(_13067_));
 sky130_fd_sc_hd__inv_1 _20153_ (.A(_11762_),
    .Y(_13071_));
 sky130_fd_sc_hd__inv_1 _20154_ (.A(_11770_),
    .Y(_13075_));
 sky130_fd_sc_hd__inv_1 _20155_ (.A(_11778_),
    .Y(_13079_));
 sky130_fd_sc_hd__inv_1 _20156_ (.A(_11786_),
    .Y(_13083_));
 sky130_fd_sc_hd__inv_2 _20157_ (.A(_11794_),
    .Y(_13087_));
 sky130_fd_sc_hd__inv_1 _20158_ (.A(_11802_),
    .Y(_13091_));
 sky130_fd_sc_hd__inv_1 _20159_ (.A(_11810_),
    .Y(_13095_));
 sky130_fd_sc_hd__clkinv_1 _20160_ (.A(_11818_),
    .Y(_13099_));
 sky130_fd_sc_hd__clkinv_1 _20161_ (.A(_11826_),
    .Y(_13103_));
 sky130_fd_sc_hd__clkinv_1 _20162_ (.A(_11831_),
    .Y(_13107_));
 sky130_fd_sc_hd__inv_1 _20163_ (.A(_11839_),
    .Y(_13110_));
 sky130_fd_sc_hd__inv_1 _20164_ (.A(_11847_),
    .Y(_13114_));
 sky130_fd_sc_hd__inv_1 _20165_ (.A(_11858_),
    .Y(_13118_));
 sky130_fd_sc_hd__inv_1 _20166_ (.A(_11866_),
    .Y(_13122_));
 sky130_fd_sc_hd__inv_1 _20167_ (.A(_11874_),
    .Y(_13126_));
 sky130_fd_sc_hd__inv_1 _20168_ (.A(_11882_),
    .Y(_13130_));
 sky130_fd_sc_hd__inv_1 _20169_ (.A(_11890_),
    .Y(_13134_));
 sky130_fd_sc_hd__inv_1 _20170_ (.A(_11898_),
    .Y(_13138_));
 sky130_fd_sc_hd__inv_1 _20171_ (.A(_11906_),
    .Y(_13142_));
 sky130_fd_sc_hd__clkinv_1 _20172_ (.A(_11914_),
    .Y(_13146_));
 sky130_fd_sc_hd__inv_1 _20173_ (.A(_11922_),
    .Y(_13150_));
 sky130_fd_sc_hd__inv_1 _20174_ (.A(_11930_),
    .Y(_13154_));
 sky130_fd_sc_hd__inv_1 _20175_ (.A(_11938_),
    .Y(_13158_));
 sky130_fd_sc_hd__inv_1 _20176_ (.A(_11946_),
    .Y(_13162_));
 sky130_fd_sc_hd__inv_1 _20177_ (.A(_11954_),
    .Y(_13166_));
 sky130_fd_sc_hd__inv_1 _20178_ (.A(_11962_),
    .Y(_13170_));
 sky130_fd_sc_hd__clkinv_1 _20179_ (.A(_11970_),
    .Y(_13174_));
 sky130_fd_sc_hd__inv_2 _20180_ (.A(_11978_),
    .Y(_13178_));
 sky130_fd_sc_hd__inv_2 _20181_ (.A(_11986_),
    .Y(_13182_));
 sky130_fd_sc_hd__inv_1 _20182_ (.A(_11994_),
    .Y(_13186_));
 sky130_fd_sc_hd__inv_1 _20183_ (.A(_12002_),
    .Y(_13190_));
 sky130_fd_sc_hd__inv_1 _20184_ (.A(_12010_),
    .Y(_13194_));
 sky130_fd_sc_hd__clkinv_1 _20185_ (.A(_12018_),
    .Y(_13198_));
 sky130_fd_sc_hd__inv_1 _20186_ (.A(_12026_),
    .Y(_13202_));
 sky130_fd_sc_hd__inv_1 _20187_ (.A(_12034_),
    .Y(_13206_));
 sky130_fd_sc_hd__inv_1 _20188_ (.A(_12042_),
    .Y(_13210_));
 sky130_fd_sc_hd__inv_1 _20189_ (.A(_12050_),
    .Y(_13214_));
 sky130_fd_sc_hd__inv_1 _20190_ (.A(_12058_),
    .Y(_13218_));
 sky130_fd_sc_hd__inv_1 _20191_ (.A(_12066_),
    .Y(_13222_));
 sky130_fd_sc_hd__inv_1 _20192_ (.A(_12074_),
    .Y(_13226_));
 sky130_fd_sc_hd__inv_1 _20193_ (.A(_12079_),
    .Y(_13233_));
 sky130_fd_sc_hd__inv_1 _20194_ (.A(_12091_),
    .Y(_12093_));
 sky130_fd_sc_hd__xnor2_4 _20195_ (.A(\hash.CA2.S1.X[8] ),
    .B(\hash.CA2.S1.X[27] ),
    .Y(_08107_));
 sky130_fd_sc_hd__xnor2_2 _20196_ (.A(_08107_),
    .B(\hash.CA2.S1.X[13] ),
    .Y(_13243_));
 sky130_fd_sc_hd__inv_1 _20197_ (.A(_12100_),
    .Y(_12102_));
 sky130_fd_sc_hd__xnor2_1 _20198_ (.A(\hash.CA2.S1.X[9] ),
    .B(\hash.CA2.S1.X[28] ),
    .Y(_08108_));
 sky130_fd_sc_hd__xnor2_1 _20199_ (.A(\hash.CA2.S1.X[14] ),
    .B(_08108_),
    .Y(_13250_));
 sky130_fd_sc_hd__inv_1 _20200_ (.A(_12114_),
    .Y(_12116_));
 sky130_fd_sc_hd__xnor2_2 _20201_ (.A(\hash.CA2.S1.X[10] ),
    .B(\hash.CA2.S1.X[29] ),
    .Y(_08109_));
 sky130_fd_sc_hd__xnor2_2 _20202_ (.A(\hash.CA2.S1.X[15] ),
    .B(_08109_),
    .Y(_13257_));
 sky130_fd_sc_hd__inv_1 _20203_ (.A(_12123_),
    .Y(_12125_));
 sky130_fd_sc_hd__xnor2_1 _20204_ (.A(\hash.CA2.S1.X[16] ),
    .B(\hash.CA2.S1.X[30] ),
    .Y(_08110_));
 sky130_fd_sc_hd__xnor2_2 _20205_ (.A(\hash.CA2.S1.X[11] ),
    .B(_08110_),
    .Y(_13264_));
 sky130_fd_sc_hd__clkinv_1 _20206_ (.A(_12132_),
    .Y(_12134_));
 sky130_fd_sc_hd__xnor2_1 _20207_ (.A(\hash.CA2.S1.X[12] ),
    .B(\hash.CA2.S1.X[17] ),
    .Y(_08111_));
 sky130_fd_sc_hd__xnor2_1 _20208_ (.A(\hash.CA2.S1.X[31] ),
    .B(_08111_),
    .Y(_13271_));
 sky130_fd_sc_hd__inv_1 _20209_ (.A(_12141_),
    .Y(_12143_));
 sky130_fd_sc_hd__xnor2_1 _20210_ (.A(\hash.CA2.S1.X[13] ),
    .B(\hash.CA2.S1.X[18] ),
    .Y(_08112_));
 sky130_fd_sc_hd__xnor2_1 _20211_ (.A(\hash.CA2.S1.X[0] ),
    .B(_08112_),
    .Y(_13278_));
 sky130_fd_sc_hd__inv_1 _20212_ (.A(_12150_),
    .Y(_12152_));
 sky130_fd_sc_hd__xnor2_1 _20213_ (.A(\hash.CA2.S1.X[14] ),
    .B(\hash.CA2.S1.X[19] ),
    .Y(_08113_));
 sky130_fd_sc_hd__xnor2_1 _20214_ (.A(net1104),
    .B(_08113_),
    .Y(_13285_));
 sky130_fd_sc_hd__inv_1 _20215_ (.A(_12159_),
    .Y(_12161_));
 sky130_fd_sc_hd__xnor2_1 _20216_ (.A(\hash.CA2.S1.X[15] ),
    .B(\hash.CA2.S1.X[20] ),
    .Y(_08114_));
 sky130_fd_sc_hd__xnor2_1 _20217_ (.A(\hash.CA2.S1.X[2] ),
    .B(_08114_),
    .Y(_13292_));
 sky130_fd_sc_hd__inv_1 _20218_ (.A(_12168_),
    .Y(_12170_));
 sky130_fd_sc_hd__xnor2_1 _20219_ (.A(\hash.CA2.S1.X[16] ),
    .B(\hash.CA2.S1.X[21] ),
    .Y(_08115_));
 sky130_fd_sc_hd__xnor2_1 _20220_ (.A(\hash.CA2.S1.X[3] ),
    .B(_08115_),
    .Y(_13299_));
 sky130_fd_sc_hd__inv_1 _20221_ (.A(_12177_),
    .Y(_12179_));
 sky130_fd_sc_hd__xnor2_1 _20222_ (.A(\hash.CA2.S1.X[17] ),
    .B(\hash.CA2.S1.X[22] ),
    .Y(_08116_));
 sky130_fd_sc_hd__xnor2_1 _20223_ (.A(\hash.CA2.S1.X[4] ),
    .B(_08116_),
    .Y(_13306_));
 sky130_fd_sc_hd__clkinv_1 _20224_ (.A(_12186_),
    .Y(_12188_));
 sky130_fd_sc_hd__xnor2_1 _20225_ (.A(\hash.CA2.S1.X[18] ),
    .B(\hash.CA2.S1.X[23] ),
    .Y(_08117_));
 sky130_fd_sc_hd__xnor2_1 _20226_ (.A(\hash.CA2.S1.X[5] ),
    .B(_08117_),
    .Y(_13313_));
 sky130_fd_sc_hd__inv_1 _20227_ (.A(_12195_),
    .Y(_12197_));
 sky130_fd_sc_hd__xnor2_1 _20228_ (.A(\hash.CA2.S1.X[19] ),
    .B(\hash.CA2.S1.X[24] ),
    .Y(_08118_));
 sky130_fd_sc_hd__xnor2_1 _20229_ (.A(net1074),
    .B(_08118_),
    .Y(_13320_));
 sky130_fd_sc_hd__inv_1 _20230_ (.A(_12204_),
    .Y(_12206_));
 sky130_fd_sc_hd__xnor2_1 _20231_ (.A(net1080),
    .B(\hash.CA2.S1.X[20] ),
    .Y(_08119_));
 sky130_fd_sc_hd__xnor2_1 _20232_ (.A(net1062),
    .B(_08119_),
    .Y(_13327_));
 sky130_fd_sc_hd__inv_1 _20233_ (.A(_12213_),
    .Y(_12215_));
 sky130_fd_sc_hd__xnor2_1 _20234_ (.A(net1115),
    .B(\hash.CA2.S1.X[21] ),
    .Y(_08120_));
 sky130_fd_sc_hd__xnor2_2 _20235_ (.A(net1087),
    .B(_08120_),
    .Y(_13334_));
 sky130_fd_sc_hd__inv_1 _20236_ (.A(_12222_),
    .Y(_12224_));
 sky130_fd_sc_hd__xnor2_1 _20237_ (.A(\hash.CA2.S1.X[9] ),
    .B(\hash.CA2.S1.X[22] ),
    .Y(_08121_));
 sky130_fd_sc_hd__xnor2_2 _20238_ (.A(\hash.CA2.S1.X[27] ),
    .B(_08121_),
    .Y(_13341_));
 sky130_fd_sc_hd__inv_1 _20239_ (.A(_12231_),
    .Y(_12233_));
 sky130_fd_sc_hd__xnor2_1 _20240_ (.A(\hash.CA2.S1.X[10] ),
    .B(\hash.CA2.S1.X[23] ),
    .Y(_08122_));
 sky130_fd_sc_hd__xnor2_1 _20241_ (.A(\hash.CA2.S1.X[28] ),
    .B(_08122_),
    .Y(_13348_));
 sky130_fd_sc_hd__inv_1 _20242_ (.A(_12240_),
    .Y(_12242_));
 sky130_fd_sc_hd__xnor2_1 _20243_ (.A(\hash.CA2.S1.X[29] ),
    .B(\hash.CA2.S1.X[24] ),
    .Y(_08123_));
 sky130_fd_sc_hd__xnor2_1 _20244_ (.A(\hash.CA2.S1.X[11] ),
    .B(_08123_),
    .Y(_13355_));
 sky130_fd_sc_hd__inv_1 _20245_ (.A(_12249_),
    .Y(_12251_));
 sky130_fd_sc_hd__xnor2_1 _20246_ (.A(\hash.CA2.S1.X[12] ),
    .B(\hash.CA2.S1.X[30] ),
    .Y(_08124_));
 sky130_fd_sc_hd__xnor2_1 _20247_ (.A(net1063),
    .B(_08124_),
    .Y(_13362_));
 sky130_fd_sc_hd__inv_1 _20248_ (.A(_12258_),
    .Y(_12260_));
 sky130_fd_sc_hd__xnor2_1 _20249_ (.A(net1086),
    .B(\hash.CA2.S1.X[13] ),
    .Y(_08125_));
 sky130_fd_sc_hd__xnor2_2 _20250_ (.A(\hash.CA2.S1.X[31] ),
    .B(_08125_),
    .Y(_13369_));
 sky130_fd_sc_hd__inv_1 _20251_ (.A(_12267_),
    .Y(_12269_));
 sky130_fd_sc_hd__xnor2_1 _20252_ (.A(net1118),
    .B(\hash.CA2.S1.X[14] ),
    .Y(_08126_));
 sky130_fd_sc_hd__xnor2_1 _20253_ (.A(\hash.CA2.S1.X[0] ),
    .B(_08126_),
    .Y(_13376_));
 sky130_fd_sc_hd__inv_1 _20254_ (.A(_12276_),
    .Y(_12278_));
 sky130_fd_sc_hd__xnor2_1 _20255_ (.A(\hash.CA2.S1.X[28] ),
    .B(\hash.CA2.S1.X[15] ),
    .Y(_08127_));
 sky130_fd_sc_hd__xnor2_1 _20256_ (.A(\hash.CA2.S1.X[1] ),
    .B(_08127_),
    .Y(_13383_));
 sky130_fd_sc_hd__inv_1 _20257_ (.A(_12285_),
    .Y(_12287_));
 sky130_fd_sc_hd__xnor2_1 _20258_ (.A(\hash.CA2.S1.X[29] ),
    .B(\hash.CA2.S1.X[16] ),
    .Y(_08128_));
 sky130_fd_sc_hd__xnor2_1 _20259_ (.A(\hash.CA2.S1.X[2] ),
    .B(_08128_),
    .Y(_13390_));
 sky130_fd_sc_hd__inv_1 _20260_ (.A(_12294_),
    .Y(_12296_));
 sky130_fd_sc_hd__xnor2_1 _20261_ (.A(\hash.CA2.S1.X[30] ),
    .B(\hash.CA2.S1.X[17] ),
    .Y(_08129_));
 sky130_fd_sc_hd__xnor2_1 _20262_ (.A(\hash.CA2.S1.X[3] ),
    .B(_08129_),
    .Y(_13397_));
 sky130_fd_sc_hd__inv_1 _20263_ (.A(_12303_),
    .Y(_12305_));
 sky130_fd_sc_hd__xnor2_2 _20264_ (.A(\hash.CA2.S1.X[4] ),
    .B(\hash.CA2.S1.X[18] ),
    .Y(_08130_));
 sky130_fd_sc_hd__xnor2_1 _20265_ (.A(\hash.CA2.S1.X[31] ),
    .B(_08130_),
    .Y(_13404_));
 sky130_fd_sc_hd__inv_1 _20266_ (.A(_12312_),
    .Y(_12314_));
 sky130_fd_sc_hd__xnor2_1 _20267_ (.A(\hash.CA2.S1.X[5] ),
    .B(\hash.CA2.S1.X[19] ),
    .Y(_08131_));
 sky130_fd_sc_hd__xnor2_1 _20268_ (.A(\hash.CA2.S1.X[0] ),
    .B(_08131_),
    .Y(_13411_));
 sky130_fd_sc_hd__inv_1 _20269_ (.A(_12321_),
    .Y(_12323_));
 sky130_fd_sc_hd__xnor2_1 _20270_ (.A(net1104),
    .B(\hash.CA2.S1.X[20] ),
    .Y(_08132_));
 sky130_fd_sc_hd__xnor2_1 _20271_ (.A(net1075),
    .B(_08132_),
    .Y(_13418_));
 sky130_fd_sc_hd__inv_1 _20272_ (.A(_12330_),
    .Y(_12332_));
 sky130_fd_sc_hd__xnor2_1 _20273_ (.A(net1119),
    .B(\hash.CA2.S1.X[21] ),
    .Y(_08133_));
 sky130_fd_sc_hd__xnor2_1 _20274_ (.A(net1080),
    .B(_08133_),
    .Y(_13425_));
 sky130_fd_sc_hd__inv_1 _20275_ (.A(_12339_),
    .Y(_12341_));
 sky130_fd_sc_hd__xnor2_1 _20276_ (.A(\hash.CA2.S1.X[3] ),
    .B(\hash.CA2.S1.X[22] ),
    .Y(_08134_));
 sky130_fd_sc_hd__xnor2_1 _20277_ (.A(\hash.CA2.S1.X[8] ),
    .B(_08134_),
    .Y(_13432_));
 sky130_fd_sc_hd__inv_1 _20278_ (.A(_12348_),
    .Y(_12350_));
 sky130_fd_sc_hd__xnor2_1 _20279_ (.A(\hash.CA2.S1.X[4] ),
    .B(\hash.CA2.S1.X[23] ),
    .Y(_08135_));
 sky130_fd_sc_hd__xnor2_1 _20280_ (.A(\hash.CA2.S1.X[9] ),
    .B(_08135_),
    .Y(_13439_));
 sky130_fd_sc_hd__inv_1 _20281_ (.A(_12357_),
    .Y(_12359_));
 sky130_fd_sc_hd__inv_1 _20282_ (.A(_12087_),
    .Y(_12363_));
 sky130_fd_sc_hd__xnor2_1 _20283_ (.A(_13427_),
    .B(_04760_),
    .Y(_13428_));
 sky130_fd_sc_hd__xor2_1 _20284_ (.A(_13441_),
    .B(_04777_),
    .X(_13442_));
 sky130_fd_sc_hd__inv_2 _20285_ (.A(\count_1[2] ),
    .Y(_13527_));
 sky130_fd_sc_hd__inv_2 _20286_ (.A(\count_2[2] ),
    .Y(_13535_));
 sky130_fd_sc_hd__xnor2_1 _20287_ (.A(_06010_),
    .B(\hash.CA1.S0.X[15] ),
    .Y(_08136_));
 sky130_fd_sc_hd__xnor2_1 _20288_ (.A(_06179_),
    .B(_08136_),
    .Y(_13552_));
 sky130_fd_sc_hd__xnor2_1 _20289_ (.A(_06016_),
    .B(_06108_),
    .Y(_08137_));
 sky130_fd_sc_hd__xnor2_4 _20290_ (.A(net1049),
    .B(_08137_),
    .Y(_13556_));
 sky130_fd_sc_hd__xnor2_1 _20291_ (.A(\hash.CA1.S0.X[6] ),
    .B(\hash.CA1.S0.X[17] ),
    .Y(_08138_));
 sky130_fd_sc_hd__xnor2_1 _20292_ (.A(_06201_),
    .B(_08138_),
    .Y(_13560_));
 sky130_fd_sc_hd__xnor2_1 _20293_ (.A(\hash.CA1.S0.X[7] ),
    .B(\hash.CA1.S0.X[18] ),
    .Y(_08139_));
 sky130_fd_sc_hd__xnor2_1 _20294_ (.A(_06211_),
    .B(_08139_),
    .Y(_13564_));
 sky130_fd_sc_hd__xnor2_1 _20295_ (.A(_06043_),
    .B(_06133_),
    .Y(_08140_));
 sky130_fd_sc_hd__xnor2_1 _20296_ (.A(_06218_),
    .B(_08140_),
    .Y(_13568_));
 sky130_fd_sc_hd__xor2_1 _20297_ (.A(\hash.CA1.S0.X[9] ),
    .B(_06148_),
    .X(_08141_));
 sky130_fd_sc_hd__xnor2_1 _20298_ (.A(_06226_),
    .B(_08141_),
    .Y(_13572_));
 sky130_fd_sc_hd__xnor2_1 _20299_ (.A(\hash.CA1.S0.X[10] ),
    .B(_06156_),
    .Y(_08142_));
 sky130_fd_sc_hd__xnor2_4 _20300_ (.A(_06234_),
    .B(_08142_),
    .Y(_13576_));
 sky130_fd_sc_hd__xnor2_1 _20301_ (.A(_06066_),
    .B(\hash.CA1.S0.X[22] ),
    .Y(_08143_));
 sky130_fd_sc_hd__xnor2_1 _20302_ (.A(_06269_),
    .B(_08143_),
    .Y(_13580_));
 sky130_fd_sc_hd__xnor2_1 _20303_ (.A(_13235_),
    .B(_06073_),
    .Y(_08144_));
 sky130_fd_sc_hd__nor2_1 _20304_ (.A(net340),
    .B(_08144_),
    .Y(_08145_));
 sky130_fd_sc_hd__xor2_1 _20305_ (.A(_06172_),
    .B(_08145_),
    .X(_13584_));
 sky130_fd_sc_hd__xor2_1 _20306_ (.A(_13241_),
    .B(_06079_),
    .X(_08146_));
 sky130_fd_sc_hd__xnor2_1 _20307_ (.A(_07935_),
    .B(_08146_),
    .Y(_08147_));
 sky130_fd_sc_hd__nor2_1 _20308_ (.A(net341),
    .B(_08147_),
    .Y(_13588_));
 sky130_fd_sc_hd__xnor2_1 _20309_ (.A(_05998_),
    .B(_06091_),
    .Y(_08148_));
 sky130_fd_sc_hd__xnor2_1 _20310_ (.A(_06212_),
    .B(_08148_),
    .Y(_08149_));
 sky130_fd_sc_hd__nand2_1 _20311_ (.A(_06002_),
    .B(_08149_),
    .Y(_13592_));
 sky130_fd_sc_hd__xnor2_1 _20312_ (.A(\hash.CA1.S0.X[3] ),
    .B(\hash.CA1.S0.X[15] ),
    .Y(_08150_));
 sky130_fd_sc_hd__xnor2_1 _20313_ (.A(_06201_),
    .B(_08150_),
    .Y(_13596_));
 sky130_fd_sc_hd__xnor2_1 _20314_ (.A(_06010_),
    .B(\hash.CA1.S0.X[16] ),
    .Y(_08151_));
 sky130_fd_sc_hd__xnor2_1 _20315_ (.A(_06211_),
    .B(_08151_),
    .Y(_13600_));
 sky130_fd_sc_hd__xnor2_1 _20316_ (.A(_06016_),
    .B(\hash.CA1.S0.X[17] ),
    .Y(_08152_));
 sky130_fd_sc_hd__xnor2_1 _20317_ (.A(_06218_),
    .B(_08152_),
    .Y(_13604_));
 sky130_fd_sc_hd__xnor2_1 _20318_ (.A(_06024_),
    .B(\hash.CA1.S0.X[18] ),
    .Y(_08153_));
 sky130_fd_sc_hd__xnor2_1 _20319_ (.A(_06226_),
    .B(_08153_),
    .Y(_13608_));
 sky130_fd_sc_hd__xnor2_1 _20320_ (.A(_06032_),
    .B(_06133_),
    .Y(_08154_));
 sky130_fd_sc_hd__xnor2_1 _20321_ (.A(_06234_),
    .B(_08154_),
    .Y(_13612_));
 sky130_fd_sc_hd__xor2_1 _20322_ (.A(_06043_),
    .B(_06148_),
    .X(_08155_));
 sky130_fd_sc_hd__xnor2_4 _20323_ (.A(_08155_),
    .B(_06269_),
    .Y(_13616_));
 sky130_fd_sc_hd__xnor2_1 _20324_ (.A(_13235_),
    .B(_06155_),
    .Y(_08156_));
 sky130_fd_sc_hd__nand2_1 _20325_ (.A(_06002_),
    .B(_08156_),
    .Y(_08157_));
 sky130_fd_sc_hd__xor2_1 _20326_ (.A(\hash.CA1.S0.X[9] ),
    .B(_08157_),
    .X(_13620_));
 sky130_fd_sc_hd__xnor2_1 _20327_ (.A(_13241_),
    .B(net1127),
    .Y(_08158_));
 sky130_fd_sc_hd__nor2_1 _20328_ (.A(net340),
    .B(_08158_),
    .Y(_08159_));
 sky130_fd_sc_hd__xnor2_1 _20329_ (.A(\hash.CA1.S0.X[10] ),
    .B(_08159_),
    .Y(_13624_));
 sky130_fd_sc_hd__nor2_1 _20330_ (.A(_12109_),
    .B(_06172_),
    .Y(_08160_));
 sky130_fd_sc_hd__a21oi_2 _20331_ (.A1(_05999_),
    .A2(_06172_),
    .B1(_08160_),
    .Y(_08161_));
 sky130_fd_sc_hd__xnor2_1 _20332_ (.A(_06066_),
    .B(_08161_),
    .Y(_13628_));
 sky130_fd_sc_hd__xnor2_1 _20333_ (.A(\hash.CA1.S0.X[3] ),
    .B(\hash.CA1.S0.X[12] ),
    .Y(_08162_));
 sky130_fd_sc_hd__xnor2_1 _20334_ (.A(_06179_),
    .B(_08162_),
    .Y(_13632_));
 sky130_fd_sc_hd__xor2_1 _20335_ (.A(_06010_),
    .B(_06080_),
    .X(_08163_));
 sky130_fd_sc_hd__xnor2_1 _20336_ (.A(net1049),
    .B(_08163_),
    .Y(_13636_));
 sky130_fd_sc_hd__xnor2_1 _20337_ (.A(\hash.CA1.S0.X[5] ),
    .B(\hash.CA1.S0.X[14] ),
    .Y(_08164_));
 sky130_fd_sc_hd__xnor2_1 _20338_ (.A(_06201_),
    .B(_08164_),
    .Y(_13640_));
 sky130_fd_sc_hd__xnor2_1 _20339_ (.A(\hash.CA1.S0.X[6] ),
    .B(\hash.CA1.S0.X[15] ),
    .Y(_08165_));
 sky130_fd_sc_hd__xnor2_1 _20340_ (.A(_06211_),
    .B(_08165_),
    .Y(_13644_));
 sky130_fd_sc_hd__xnor2_1 _20341_ (.A(\hash.CA1.S0.X[7] ),
    .B(_06108_),
    .Y(_08166_));
 sky130_fd_sc_hd__xnor2_1 _20342_ (.A(_06218_),
    .B(_08166_),
    .Y(_13648_));
 sky130_fd_sc_hd__xor2_1 _20343_ (.A(_06043_),
    .B(\hash.CA1.S0.X[17] ),
    .X(_08167_));
 sky130_fd_sc_hd__xnor2_1 _20344_ (.A(_06226_),
    .B(_08167_),
    .Y(_13652_));
 sky130_fd_sc_hd__xnor2_1 _20345_ (.A(\hash.CA1.S0.X[9] ),
    .B(\hash.CA1.S0.X[18] ),
    .Y(_08168_));
 sky130_fd_sc_hd__xnor2_1 _20346_ (.A(_06234_),
    .B(_08168_),
    .Y(_13656_));
 sky130_fd_sc_hd__xnor2_1 _20347_ (.A(\hash.CA1.S0.X[10] ),
    .B(_06133_),
    .Y(_08169_));
 sky130_fd_sc_hd__xnor2_1 _20348_ (.A(_06269_),
    .B(_08169_),
    .Y(_13660_));
 sky130_fd_sc_hd__mux2i_1 _20349_ (.A0(_13235_),
    .A1(_00658_),
    .S(_06066_),
    .Y(_08170_));
 sky130_fd_sc_hd__xor2_1 _20350_ (.A(_06148_),
    .B(_08170_),
    .X(_13664_));
 sky130_fd_sc_hd__inv_1 _20351_ (.A(_12370_),
    .Y(_13668_));
 sky130_fd_sc_hd__inv_1 _20352_ (.A(_12385_),
    .Y(_13676_));
 sky130_fd_sc_hd__inv_1 _20353_ (.A(_12393_),
    .Y(_13688_));
 sky130_fd_sc_hd__inv_1 _20354_ (.A(_12401_),
    .Y(_13700_));
 sky130_fd_sc_hd__inv_1 _20355_ (.A(_06800_),
    .Y(_13703_));
 sky130_fd_sc_hd__inv_1 _20356_ (.A(_12406_),
    .Y(_13707_));
 sky130_fd_sc_hd__clkinv_1 _20357_ (.A(_12417_),
    .Y(_13724_));
 sky130_fd_sc_hd__nor2b_1 _20358_ (.A(net346),
    .B_N(\hash.CA2.a_dash[11] ),
    .Y(_13727_));
 sky130_fd_sc_hd__inv_1 _20359_ (.A(_12422_),
    .Y(_13731_));
 sky130_fd_sc_hd__inv_1 _20360_ (.A(_12430_),
    .Y(_13743_));
 sky130_fd_sc_hd__inv_1 _20361_ (.A(_12435_),
    .Y(_13750_));
 sky130_fd_sc_hd__inv_1 _20362_ (.A(_12440_),
    .Y(_13757_));
 sky130_fd_sc_hd__inv_1 _20363_ (.A(_12445_),
    .Y(_13764_));
 sky130_fd_sc_hd__inv_1 _20364_ (.A(_12465_),
    .Y(_13796_));
 sky130_fd_sc_hd__inv_1 _20365_ (.A(_12470_),
    .Y(_13803_));
 sky130_fd_sc_hd__nor2b_1 _20366_ (.A(net346),
    .B_N(\hash.CA2.a_dash[24] ),
    .Y(_13806_));
 sky130_fd_sc_hd__inv_1 _20367_ (.A(_12475_),
    .Y(_13810_));
 sky130_fd_sc_hd__nor2_1 _20368_ (.A(net346),
    .B(_04734_),
    .Y(_13813_));
 sky130_fd_sc_hd__inv_1 _20369_ (.A(_12480_),
    .Y(_13817_));
 sky130_fd_sc_hd__inv_1 _20370_ (.A(_12485_),
    .Y(_13824_));
 sky130_fd_sc_hd__inv_1 _20371_ (.A(_12490_),
    .Y(_13831_));
 sky130_fd_sc_hd__mux2i_2 _20372_ (.A0(\hash.CA2.e_dash[2] ),
    .A1(\hash.CA2.S1.X[2] ),
    .S(_06513_),
    .Y(_08171_));
 sky130_fd_sc_hd__nand2_2 _20373_ (.A(_06002_),
    .B(_08171_),
    .Y(_13870_));
 sky130_fd_sc_hd__inv_1 _20374_ (.A(_12517_),
    .Y(_13881_));
 sky130_fd_sc_hd__mux2_8 _20375_ (.A0(\hash.CA1.f[4] ),
    .A1(\hash.CA2.e_dash[4] ),
    .S(_06524_),
    .X(_13887_));
 sky130_fd_sc_hd__inv_1 _20376_ (.A(_12522_),
    .Y(_13891_));
 sky130_fd_sc_hd__nand2_1 _20377_ (.A(\hash.CA2.e_dash[5] ),
    .B(_06531_),
    .Y(_08172_));
 sky130_fd_sc_hd__nand2_1 _20378_ (.A(\hash.CA1.f[5] ),
    .B(\hash.CA1.S1.X[5] ),
    .Y(_08173_));
 sky130_fd_sc_hd__nand2_4 _20379_ (.A(_08172_),
    .B(_08173_),
    .Y(_13897_));
 sky130_fd_sc_hd__mux2i_4 _20380_ (.A0(_12399_),
    .A1(_06428_),
    .S(\hash.CA1.S1.X[7] ),
    .Y(_13914_));
 sky130_fd_sc_hd__nor3_2 _20381_ (.A(net344),
    .B(\hash.CA2.e_dash[8] ),
    .C(_06551_),
    .Y(_08174_));
 sky130_fd_sc_hd__a21oi_4 _20382_ (.A1(_06433_),
    .A2(_06552_),
    .B1(_08174_),
    .Y(_13922_));
 sky130_fd_sc_hd__inv_1 _20383_ (.A(_12542_),
    .Y(_13925_));
 sky130_fd_sc_hd__nand2_2 _20384_ (.A(\hash.CA2.e_dash[9] ),
    .B(_06559_),
    .Y(_08175_));
 sky130_fd_sc_hd__nand2_1 _20385_ (.A(_06438_),
    .B(\hash.CA1.S1.X[9] ),
    .Y(_08176_));
 sky130_fd_sc_hd__nand2_2 _20386_ (.A(_08175_),
    .B(_08176_),
    .Y(_13931_));
 sky130_fd_sc_hd__nand2_1 _20387_ (.A(\hash.CA2.S1.X[10] ),
    .B(\hash.CA1.S1.X[10] ),
    .Y(_08177_));
 sky130_fd_sc_hd__nand2_2 _20388_ (.A(_12410_),
    .B(_06568_),
    .Y(_08178_));
 sky130_fd_sc_hd__nand2_2 _20389_ (.A(_08177_),
    .B(_08178_),
    .Y(_13940_));
 sky130_fd_sc_hd__inv_2 _20390_ (.A(_12552_),
    .Y(_13943_));
 sky130_fd_sc_hd__inv_1 _20391_ (.A(_12557_),
    .Y(_13953_));
 sky130_fd_sc_hd__nand2_1 _20392_ (.A(\hash.CA2.e_dash[12] ),
    .B(_06581_),
    .Y(_08179_));
 sky130_fd_sc_hd__nand2_1 _20393_ (.A(\hash.CA1.f[12] ),
    .B(\hash.CA1.S1.X[12] ),
    .Y(_08180_));
 sky130_fd_sc_hd__nand2_1 _20394_ (.A(_08179_),
    .B(_08180_),
    .Y(_13959_));
 sky130_fd_sc_hd__nand2_2 _20395_ (.A(\hash.CA2.S1.X[13] ),
    .B(\hash.CA1.S1.X[13] ),
    .Y(_08181_));
 sky130_fd_sc_hd__nand2_4 _20396_ (.A(_12423_),
    .B(_06589_),
    .Y(_08182_));
 sky130_fd_sc_hd__nand2_4 _20397_ (.A(_08181_),
    .B(_08182_),
    .Y(_13968_));
 sky130_fd_sc_hd__inv_2 _20398_ (.A(_12572_),
    .Y(_13979_));
 sky130_fd_sc_hd__inv_1 _20399_ (.A(\hash.CA2.S1.X[15] ),
    .Y(_08183_));
 sky130_fd_sc_hd__nor3_2 _20400_ (.A(net534),
    .B(\hash.CA2.e_dash[15] ),
    .C(_06610_),
    .Y(_08184_));
 sky130_fd_sc_hd__a21oi_4 _20401_ (.A1(_08183_),
    .A2(_06610_),
    .B1(_08184_),
    .Y(_13985_));
 sky130_fd_sc_hd__inv_1 _20402_ (.A(_12577_),
    .Y(_13989_));
 sky130_fd_sc_hd__mux2_8 _20403_ (.A0(\hash.CA1.f[17] ),
    .A1(\hash.CA2.e_dash[17] ),
    .S(_06624_),
    .X(_14004_));
 sky130_fd_sc_hd__mux2_8 _20404_ (.A0(\hash.CA1.f[19] ),
    .A1(\hash.CA2.e_dash[19] ),
    .S(_06642_),
    .X(_14020_));
 sky130_fd_sc_hd__mux2_4 _20405_ (.A0(_12452_),
    .A1(\hash.CA2.S1.X[20] ),
    .S(\hash.CA1.S1.X[20] ),
    .X(_14028_));
 sky130_fd_sc_hd__mux2_4 _20406_ (.A0(_12455_),
    .A1(\hash.CA2.S1.X[21] ),
    .S(\hash.CA1.S1.X[21] ),
    .X(_14036_));
 sky130_fd_sc_hd__inv_1 _20407_ (.A(_12607_),
    .Y(_14039_));
 sky130_fd_sc_hd__mux2_1 _20408_ (.A0(_12458_),
    .A1(\hash.CA2.S1.X[22] ),
    .S(\hash.CA1.S1.X[22] ),
    .X(_14045_));
 sky130_fd_sc_hd__inv_1 _20409_ (.A(_12612_),
    .Y(_14049_));
 sky130_fd_sc_hd__nor2_1 _20410_ (.A(\hash.CA2.S1.X[23] ),
    .B(_06665_),
    .Y(_08185_));
 sky130_fd_sc_hd__a21oi_1 _20411_ (.A1(_12463_),
    .A2(_06665_),
    .B1(_08185_),
    .Y(_14055_));
 sky130_fd_sc_hd__inv_2 _20412_ (.A(_12617_),
    .Y(_14059_));
 sky130_fd_sc_hd__inv_2 _20413_ (.A(_12622_),
    .Y(_14069_));
 sky130_fd_sc_hd__inv_1 _20414_ (.A(_12627_),
    .Y(_14079_));
 sky130_fd_sc_hd__clkinvlp_2 _20415_ (.A(net1086),
    .Y(_08186_));
 sky130_fd_sc_hd__nor3_1 _20416_ (.A(net534),
    .B(\hash.CA2.e_dash[26] ),
    .C(net1056),
    .Y(_08187_));
 sky130_fd_sc_hd__a21oi_4 _20417_ (.A1(_08186_),
    .A2(net1058),
    .B1(_08187_),
    .Y(_14085_));
 sky130_fd_sc_hd__inv_1 _20418_ (.A(_12637_),
    .Y(_14097_));
 sky130_fd_sc_hd__inv_1 _20419_ (.A(_12642_),
    .Y(_14107_));
 sky130_fd_sc_hd__mux2_8 _20420_ (.A0(\hash.CA2.S1.X[29] ),
    .A1(_12491_),
    .S(_06712_),
    .X(_14113_));
 sky130_fd_sc_hd__mux2_8 _20421_ (.A0(\hash.CA2.e_dash[30] ),
    .A1(\hash.CA1.f[30] ),
    .S(net1042),
    .X(_14122_));
 sky130_fd_sc_hd__inv_1 _20422_ (.A(_12652_),
    .Y(_14125_));
 sky130_fd_sc_hd__inv_1 _20423_ (.A(_12673_),
    .Y(_14129_));
 sky130_fd_sc_hd__inv_1 _20424_ (.A(_12678_),
    .Y(_14133_));
 sky130_fd_sc_hd__inv_1 _20425_ (.A(_12683_),
    .Y(_14137_));
 sky130_fd_sc_hd__clkinv_1 _20426_ (.A(_12690_),
    .Y(_14141_));
 sky130_fd_sc_hd__clkinv_1 _20427_ (.A(_12699_),
    .Y(_14145_));
 sky130_fd_sc_hd__inv_2 _20428_ (.A(_12707_),
    .Y(_14149_));
 sky130_fd_sc_hd__inv_1 _20429_ (.A(_12712_),
    .Y(_14153_));
 sky130_fd_sc_hd__inv_1 _20430_ (.A(_12717_),
    .Y(_12719_));
 sky130_fd_sc_hd__inv_1 _20431_ (.A(_12754_),
    .Y(_12755_));
 sky130_fd_sc_hd__inv_1 _20432_ (.A(_12761_),
    .Y(_12763_));
 sky130_fd_sc_hd__inv_1 _20433_ (.A(_12796_),
    .Y(_12797_));
 sky130_fd_sc_hd__inv_1 _20434_ (.A(_12812_),
    .Y(_12813_));
 sky130_fd_sc_hd__inv_1 _20435_ (.A(_12828_),
    .Y(_12829_));
 sky130_fd_sc_hd__inv_1 _20436_ (.A(_12878_),
    .Y(_14199_));
 sky130_fd_sc_hd__xnor2_1 _20437_ (.A(_05998_),
    .B(_06079_),
    .Y(_08188_));
 sky130_fd_sc_hd__xnor2_1 _20438_ (.A(net1127),
    .B(_08188_),
    .Y(_08189_));
 sky130_fd_sc_hd__nor2_1 _20439_ (.A(net340),
    .B(_08189_),
    .Y(_14203_));
 sky130_fd_sc_hd__inv_1 _20440_ (.A(_12664_),
    .Y(_14206_));
 sky130_fd_sc_hd__inv_1 _20441_ (.A(_12374_),
    .Y(\hash.CA1.p4[0] ));
 sky130_fd_sc_hd__inv_6 _20442_ (.A(_13232_),
    .Y(_12076_));
 sky130_fd_sc_hd__inv_1 _20443_ (.A(_13856_),
    .Y(_00792_));
 sky130_fd_sc_hd__inv_1 _20444_ (.A(_13545_),
    .Y(_00669_));
 sky130_fd_sc_hd__inv_1 _20445_ (.A(\hash.CA1.p4[1] ),
    .Y(_12895_));
 sky130_fd_sc_hd__inv_1 _20446_ (.A(_13850_),
    .Y(_00854_));
 sky130_fd_sc_hd__inv_1 _20447_ (.A(_13853_),
    .Y(_00824_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_983 ();
 sky130_fd_sc_hd__nor2_1 _20449_ (.A(net1038),
    .B(net532),
    .Y(_00907_));
 sky130_fd_sc_hd__nor2b_1 _20450_ (.A(net1038),
    .B_N(_00644_),
    .Y(_00908_));
 sky130_fd_sc_hd__xnor2_1 _20451_ (.A(net518),
    .B(_13521_),
    .Y(_08191_));
 sky130_fd_sc_hd__nor2_1 _20452_ (.A(net1038),
    .B(_08191_),
    .Y(_00909_));
 sky130_fd_sc_hd__nand3_1 _20453_ (.A(net550),
    .B(\count15_1[2] ),
    .C(net518),
    .Y(_08192_));
 sky130_fd_sc_hd__xor2_1 _20454_ (.A(net549),
    .B(_08192_),
    .X(_08193_));
 sky130_fd_sc_hd__nor2_1 _20455_ (.A(net1038),
    .B(_08193_),
    .Y(_00910_));
 sky130_fd_sc_hd__nand3_1 _20456_ (.A(net518),
    .B(net515),
    .C(_13521_),
    .Y(_08194_));
 sky130_fd_sc_hd__xor2_1 _20457_ (.A(net513),
    .B(_08194_),
    .X(_08195_));
 sky130_fd_sc_hd__nor2_1 _20458_ (.A(net1038),
    .B(_08195_),
    .Y(_00911_));
 sky130_fd_sc_hd__nand2_1 _20459_ (.A(_09731_),
    .B(\count15_2[1] ),
    .Y(_00912_));
 sky130_fd_sc_hd__nor2b_1 _20460_ (.A(net780),
    .B_N(_00648_),
    .Y(_00913_));
 sky130_fd_sc_hd__xnor2_1 _20461_ (.A(\count15_2[3] ),
    .B(_13525_),
    .Y(_08196_));
 sky130_fd_sc_hd__nor2_1 _20462_ (.A(net1039),
    .B(_08196_),
    .Y(_00914_));
 sky130_fd_sc_hd__nand3_1 _20463_ (.A(\count15_2[1] ),
    .B(net505),
    .C(net497),
    .Y(_08197_));
 sky130_fd_sc_hd__xor2_1 _20464_ (.A(\count15_2[4] ),
    .B(_08197_),
    .X(_08198_));
 sky130_fd_sc_hd__nor2_1 _20465_ (.A(net1038),
    .B(_08198_),
    .Y(_00915_));
 sky130_fd_sc_hd__nand3_1 _20466_ (.A(\count15_2[3] ),
    .B(\count15_2[4] ),
    .C(_13525_),
    .Y(_08199_));
 sky130_fd_sc_hd__xor2_1 _20467_ (.A(\count15_2[5] ),
    .B(_08199_),
    .X(_08200_));
 sky130_fd_sc_hd__nor2_1 _20468_ (.A(net1039),
    .B(_08200_),
    .Y(_00916_));
 sky130_fd_sc_hd__nor2_1 _20469_ (.A(net780),
    .B(\count16_1[1] ),
    .Y(_00917_));
 sky130_fd_sc_hd__nor2b_1 _20470_ (.A(net1038),
    .B_N(_00645_),
    .Y(_00918_));
 sky130_fd_sc_hd__xnor2_1 _20471_ (.A(\count16_1[3] ),
    .B(_13522_),
    .Y(_08201_));
 sky130_fd_sc_hd__nor2_1 _20472_ (.A(net1038),
    .B(_08201_),
    .Y(_00919_));
 sky130_fd_sc_hd__nand3_1 _20473_ (.A(net490),
    .B(net484),
    .C(net477),
    .Y(_08202_));
 sky130_fd_sc_hd__xor2_1 _20474_ (.A(\count16_1[4] ),
    .B(_08202_),
    .X(_08203_));
 sky130_fd_sc_hd__nor2_1 _20475_ (.A(net1038),
    .B(_08203_),
    .Y(_00920_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_982 ();
 sky130_fd_sc_hd__nand3_1 _20477_ (.A(\count16_1[3] ),
    .B(\count16_1[4] ),
    .C(_13522_),
    .Y(_08205_));
 sky130_fd_sc_hd__xor2_1 _20478_ (.A(\count16_1[5] ),
    .B(_08205_),
    .X(_08206_));
 sky130_fd_sc_hd__nor2_1 _20479_ (.A(net1038),
    .B(_08206_),
    .Y(_00921_));
 sky130_fd_sc_hd__nor2_1 _20480_ (.A(net780),
    .B(\count16_2[1] ),
    .Y(_00922_));
 sky130_fd_sc_hd__nor2b_1 _20481_ (.A(net1038),
    .B_N(_00649_),
    .Y(_00923_));
 sky130_fd_sc_hd__xnor2_1 _20482_ (.A(net457),
    .B(_13526_),
    .Y(_08207_));
 sky130_fd_sc_hd__nor2_1 _20483_ (.A(net1038),
    .B(_08207_),
    .Y(_00924_));
 sky130_fd_sc_hd__nand3_1 _20484_ (.A(net471),
    .B(net466),
    .C(net457),
    .Y(_08208_));
 sky130_fd_sc_hd__xor2_1 _20485_ (.A(\count16_2[4] ),
    .B(_08208_),
    .X(_08209_));
 sky130_fd_sc_hd__nor2_1 _20486_ (.A(net1038),
    .B(_08209_),
    .Y(_00925_));
 sky130_fd_sc_hd__nand3_1 _20487_ (.A(\count16_2[3] ),
    .B(net455),
    .C(_13526_),
    .Y(_08210_));
 sky130_fd_sc_hd__xor2_1 _20488_ (.A(\count16_2[5] ),
    .B(_08210_),
    .X(_08211_));
 sky130_fd_sc_hd__nor2_1 _20489_ (.A(net1038),
    .B(_08211_),
    .Y(_00926_));
 sky130_fd_sc_hd__nand2_1 _20490_ (.A(_09731_),
    .B(\count2_1[1] ),
    .Y(_00927_));
 sky130_fd_sc_hd__or2_0 _20491_ (.A(net1038),
    .B(_00642_),
    .X(_00928_));
 sky130_fd_sc_hd__xnor2_1 _20492_ (.A(\count2_1[3] ),
    .B(_13546_),
    .Y(_08212_));
 sky130_fd_sc_hd__nand2_1 _20493_ (.A(_09731_),
    .B(_08212_),
    .Y(_00929_));
 sky130_fd_sc_hd__nand3_1 _20494_ (.A(net452),
    .B(\count2_1[2] ),
    .C(net438),
    .Y(_08213_));
 sky130_fd_sc_hd__xor2_1 _20495_ (.A(\count2_1[4] ),
    .B(_08213_),
    .X(_08214_));
 sky130_fd_sc_hd__nor2_1 _20496_ (.A(net1038),
    .B(_08214_),
    .Y(_00930_));
 sky130_fd_sc_hd__nand3_1 _20497_ (.A(\count2_1[3] ),
    .B(\count2_1[4] ),
    .C(_13546_),
    .Y(_08215_));
 sky130_fd_sc_hd__xor2_1 _20498_ (.A(\count2_1[5] ),
    .B(_08215_),
    .X(_08216_));
 sky130_fd_sc_hd__nor2_1 _20499_ (.A(net1038),
    .B(_08216_),
    .Y(_00931_));
 sky130_fd_sc_hd__nand2_1 _20500_ (.A(_09731_),
    .B(\count2_2[1] ),
    .Y(_00932_));
 sky130_fd_sc_hd__or2_0 _20501_ (.A(net1039),
    .B(_00646_),
    .X(_00933_));
 sky130_fd_sc_hd__xnor2_1 _20502_ (.A(\count2_2[3] ),
    .B(_13523_),
    .Y(_08217_));
 sky130_fd_sc_hd__nand2_1 _20503_ (.A(_09731_),
    .B(_08217_),
    .Y(_00934_));
 sky130_fd_sc_hd__nand3_1 _20504_ (.A(net430),
    .B(net425),
    .C(net418),
    .Y(_08218_));
 sky130_fd_sc_hd__xor2_1 _20505_ (.A(\count2_2[4] ),
    .B(_08218_),
    .X(_08219_));
 sky130_fd_sc_hd__nor2_1 _20506_ (.A(net1038),
    .B(_08219_),
    .Y(_00935_));
 sky130_fd_sc_hd__nand3_1 _20507_ (.A(\count2_2[3] ),
    .B(\count2_2[4] ),
    .C(_13523_),
    .Y(_08220_));
 sky130_fd_sc_hd__xor2_1 _20508_ (.A(\count2_2[5] ),
    .B(_08220_),
    .X(_08221_));
 sky130_fd_sc_hd__nor2_1 _20509_ (.A(net1039),
    .B(_08221_),
    .Y(_00936_));
 sky130_fd_sc_hd__nor2_1 _20510_ (.A(net780),
    .B(\count7_1[1] ),
    .Y(_00937_));
 sky130_fd_sc_hd__nor2b_1 _20511_ (.A(net1038),
    .B_N(_00643_),
    .Y(_00938_));
 sky130_fd_sc_hd__xnor2_1 _20512_ (.A(net400),
    .B(_13520_),
    .Y(_08222_));
 sky130_fd_sc_hd__nand2_1 _20513_ (.A(_09731_),
    .B(_08222_),
    .Y(_00939_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_981 ();
 sky130_fd_sc_hd__nand3_1 _20515_ (.A(net412),
    .B(\count7_1[2] ),
    .C(net537),
    .Y(_08224_));
 sky130_fd_sc_hd__xor2_1 _20516_ (.A(\count7_1[4] ),
    .B(_08224_),
    .X(_08225_));
 sky130_fd_sc_hd__nor2_1 _20517_ (.A(net1038),
    .B(_08225_),
    .Y(_00940_));
 sky130_fd_sc_hd__nand3_2 _20518_ (.A(net400),
    .B(\count7_1[4] ),
    .C(_13520_),
    .Y(_08226_));
 sky130_fd_sc_hd__xor2_1 _20519_ (.A(\count7_1[5] ),
    .B(_08226_),
    .X(_08227_));
 sky130_fd_sc_hd__nor2_1 _20520_ (.A(net1038),
    .B(_08227_),
    .Y(_00941_));
 sky130_fd_sc_hd__nand2_1 _20521_ (.A(_09731_),
    .B(\count7_2[1] ),
    .Y(_00942_));
 sky130_fd_sc_hd__nor2b_1 _20522_ (.A(net1038),
    .B_N(_00647_),
    .Y(_00943_));
 sky130_fd_sc_hd__xnor2_1 _20523_ (.A(\count7_2[3] ),
    .B(_13524_),
    .Y(_08228_));
 sky130_fd_sc_hd__nand2_1 _20524_ (.A(_09731_),
    .B(_08228_),
    .Y(_00944_));
 sky130_fd_sc_hd__nand3_1 _20525_ (.A(net393),
    .B(\count7_2[2] ),
    .C(net378),
    .Y(_08229_));
 sky130_fd_sc_hd__xor2_1 _20526_ (.A(net376),
    .B(_08229_),
    .X(_08230_));
 sky130_fd_sc_hd__nor2_1 _20527_ (.A(net1038),
    .B(_08230_),
    .Y(_00945_));
 sky130_fd_sc_hd__nand3_1 _20528_ (.A(\count7_2[3] ),
    .B(net376),
    .C(_13524_),
    .Y(_08231_));
 sky130_fd_sc_hd__xor2_1 _20529_ (.A(\count7_2[5] ),
    .B(_08231_),
    .X(_08232_));
 sky130_fd_sc_hd__nor2_1 _20530_ (.A(net1038),
    .B(_08232_),
    .Y(_00946_));
 sky130_fd_sc_hd__xnor2_1 _20531_ (.A(_00650_),
    .B(_00128_),
    .Y(_08233_));
 sky130_fd_sc_hd__nor2_1 _20532_ (.A(net780),
    .B(_08233_),
    .Y(_00947_));
 sky130_fd_sc_hd__nand2_1 _20533_ (.A(\count_1[2] ),
    .B(_00128_),
    .Y(_08234_));
 sky130_fd_sc_hd__nand2_1 _20534_ (.A(_00651_),
    .B(_09727_),
    .Y(_08235_));
 sky130_fd_sc_hd__a21oi_1 _20535_ (.A1(_08234_),
    .A2(_08235_),
    .B1(net780),
    .Y(_00948_));
 sky130_fd_sc_hd__nand2_1 _20536_ (.A(_13533_),
    .B(_09727_),
    .Y(_08236_));
 sky130_fd_sc_hd__xor2_1 _20537_ (.A(\count_1[3] ),
    .B(_08236_),
    .X(_08237_));
 sky130_fd_sc_hd__nor2_1 _20538_ (.A(net1039),
    .B(_08237_),
    .Y(_00949_));
 sky130_fd_sc_hd__nand4_1 _20539_ (.A(\count_1[3] ),
    .B(\count_1[2] ),
    .C(\count_1[1] ),
    .D(_09727_),
    .Y(_08238_));
 sky130_fd_sc_hd__xor2_1 _20540_ (.A(\count_1[4] ),
    .B(_08238_),
    .X(_08239_));
 sky130_fd_sc_hd__nand2_1 _20541_ (.A(_09731_),
    .B(_08239_),
    .Y(_00950_));
 sky130_fd_sc_hd__nand4_1 _20542_ (.A(\count_1[4] ),
    .B(\count_1[3] ),
    .C(_13533_),
    .D(_09727_),
    .Y(_08240_));
 sky130_fd_sc_hd__xor2_1 _20543_ (.A(\count_1[5] ),
    .B(_08240_),
    .X(_08241_));
 sky130_fd_sc_hd__nor2_1 _20544_ (.A(net1039),
    .B(_08241_),
    .Y(_00951_));
 sky130_fd_sc_hd__xnor2_1 _20545_ (.A(_00652_),
    .B(_00128_),
    .Y(_08242_));
 sky130_fd_sc_hd__nor2_1 _20546_ (.A(net1039),
    .B(_08242_),
    .Y(_00952_));
 sky130_fd_sc_hd__nand2_1 _20547_ (.A(\count_2[2] ),
    .B(_00128_),
    .Y(_08243_));
 sky130_fd_sc_hd__nand2_1 _20548_ (.A(_00653_),
    .B(_09727_),
    .Y(_08244_));
 sky130_fd_sc_hd__a21oi_1 _20549_ (.A1(_08243_),
    .A2(_08244_),
    .B1(net1039),
    .Y(_00953_));
 sky130_fd_sc_hd__xnor2_1 _20550_ (.A(\count_2[3] ),
    .B(_13541_),
    .Y(_08245_));
 sky130_fd_sc_hd__a21oi_1 _20551_ (.A1(_09727_),
    .A2(_08245_),
    .B1(net1039),
    .Y(_00954_));
 sky130_fd_sc_hd__nand3_1 _20552_ (.A(\count_2[3] ),
    .B(\count_2[2] ),
    .C(\count_2[1] ),
    .Y(_08246_));
 sky130_fd_sc_hd__xor2_1 _20553_ (.A(\count_2[4] ),
    .B(_08246_),
    .X(_08247_));
 sky130_fd_sc_hd__nand3_1 _20554_ (.A(_09731_),
    .B(_09727_),
    .C(_08247_),
    .Y(_00955_));
 sky130_fd_sc_hd__nand3_1 _20555_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(_13541_),
    .Y(_08248_));
 sky130_fd_sc_hd__nand2_1 _20556_ (.A(\count_2[6] ),
    .B(\count_2[5] ),
    .Y(_08249_));
 sky130_fd_sc_hd__nor2_1 _20557_ (.A(_08248_),
    .B(_08249_),
    .Y(_08250_));
 sky130_fd_sc_hd__a211oi_1 _20558_ (.A1(_09802_),
    .A2(_08248_),
    .B1(_08250_),
    .C1(net1038),
    .Y(_00956_));
 sky130_fd_sc_hd__nor2b_1 _20559_ (.A(\count_2[6] ),
    .B_N(_09726_),
    .Y(_08251_));
 sky130_fd_sc_hd__nand2_1 _20560_ (.A(\count_2[4] ),
    .B(\count_2[5] ),
    .Y(_08252_));
 sky130_fd_sc_hd__nor2_1 _20561_ (.A(_08246_),
    .B(_08252_),
    .Y(_08253_));
 sky130_fd_sc_hd__mux2i_1 _20562_ (.A0(\count_2[6] ),
    .A1(_08251_),
    .S(_08253_),
    .Y(_08254_));
 sky130_fd_sc_hd__nor2_1 _20563_ (.A(net1039),
    .B(_08254_),
    .Y(_00957_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_980 ();
 sky130_fd_sc_hd__nand3_2 _20565_ (.A(\count_hash1[4] ),
    .B(\count_hash1[3] ),
    .C(\count_hash1[5] ),
    .Y(_08256_));
 sky130_fd_sc_hd__nor2_4 _20566_ (.A(\count_hash1[6] ),
    .B(_08256_),
    .Y(_08257_));
 sky130_fd_sc_hd__nand2_8 _20567_ (.A(_12920_),
    .B(_08257_),
    .Y(_08258_));
 sky130_fd_sc_hd__xnor2_1 _20568_ (.A(net372),
    .B(_08258_),
    .Y(_08259_));
 sky130_fd_sc_hd__nor2_1 _20569_ (.A(net349),
    .B(_08259_),
    .Y(_00958_));
 sky130_fd_sc_hd__nor2_1 _20570_ (.A(_12910_),
    .B(_08258_),
    .Y(_08260_));
 sky130_fd_sc_hd__a21oi_1 _20571_ (.A1(_00655_),
    .A2(_08258_),
    .B1(_08260_),
    .Y(_08261_));
 sky130_fd_sc_hd__nor2_1 _20572_ (.A(net348),
    .B(_08261_),
    .Y(_00959_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_978 ();
 sky130_fd_sc_hd__nor2_1 _20575_ (.A(net325),
    .B(_08257_),
    .Y(_08264_));
 sky130_fd_sc_hd__nor2_1 _20576_ (.A(net349),
    .B(_08264_),
    .Y(_00960_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_977 ();
 sky130_fd_sc_hd__a21oi_1 _20578_ (.A1(_10352_),
    .A2(_08258_),
    .B1(net349),
    .Y(_00961_));
 sky130_fd_sc_hd__xor2_4 _20579_ (.A(\count_hash1[5] ),
    .B(_10372_),
    .X(_08266_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_974 ();
 sky130_fd_sc_hd__a21oi_1 _20583_ (.A1(_08266_),
    .A2(_08258_),
    .B1(net349),
    .Y(_00962_));
 sky130_fd_sc_hd__or4_1 _20584_ (.A(_12920_),
    .B(_00654_),
    .C(\count_hash1[6] ),
    .D(_09873_),
    .X(_08270_));
 sky130_fd_sc_hd__o21ai_0 _20585_ (.A1(_00654_),
    .A2(_09873_),
    .B1(\count_hash1[6] ),
    .Y(_08271_));
 sky130_fd_sc_hd__a21oi_1 _20586_ (.A1(_08270_),
    .A2(_08271_),
    .B1(net349),
    .Y(_00963_));
 sky130_fd_sc_hd__xnor2_1 _20587_ (.A(\count_hash2[1] ),
    .B(_08258_),
    .Y(_08272_));
 sky130_fd_sc_hd__nor2_1 _20588_ (.A(net349),
    .B(_08272_),
    .Y(_00964_));
 sky130_fd_sc_hd__nor2_1 _20589_ (.A(_12900_),
    .B(_08258_),
    .Y(_08273_));
 sky130_fd_sc_hd__a21oi_1 _20590_ (.A1(_00657_),
    .A2(_08258_),
    .B1(_08273_),
    .Y(_08274_));
 sky130_fd_sc_hd__nor2_1 _20591_ (.A(net349),
    .B(_08274_),
    .Y(_00965_));
 sky130_fd_sc_hd__nand2_1 _20592_ (.A(_12908_),
    .B(_08258_),
    .Y(_08275_));
 sky130_fd_sc_hd__xor2_1 _20593_ (.A(\count_hash2[3] ),
    .B(_08275_),
    .X(_08276_));
 sky130_fd_sc_hd__nor2_1 _20594_ (.A(net349),
    .B(_08276_),
    .Y(_00966_));
 sky130_fd_sc_hd__a21oi_1 _20595_ (.A1(_12920_),
    .A2(_08257_),
    .B1(_09856_),
    .Y(_08277_));
 sky130_fd_sc_hd__xnor2_1 _20596_ (.A(\count_hash2[4] ),
    .B(_08277_),
    .Y(_08278_));
 sky130_fd_sc_hd__nor2_1 _20597_ (.A(net349),
    .B(_08278_),
    .Y(_00967_));
 sky130_fd_sc_hd__a21oi_1 _20598_ (.A1(_12920_),
    .A2(_08257_),
    .B1(_09866_),
    .Y(_08279_));
 sky130_fd_sc_hd__xnor2_1 _20599_ (.A(\count_hash2[5] ),
    .B(_08279_),
    .Y(_08280_));
 sky130_fd_sc_hd__nor2_1 _20600_ (.A(net349),
    .B(_08280_),
    .Y(_00968_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_972 ();
 sky130_fd_sc_hd__xnor2_4 _20603_ (.A(\count_hash1[3] ),
    .B(_12920_),
    .Y(_08283_));
 sky130_fd_sc_hd__nand2_4 _20604_ (.A(net316),
    .B(_08283_),
    .Y(_08284_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_969 ();
 sky130_fd_sc_hd__nor2_1 _20608_ (.A(_12912_),
    .B(net318),
    .Y(_08288_));
 sky130_fd_sc_hd__nor2_1 _20609_ (.A(net320),
    .B(_08288_),
    .Y(_08289_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_965 ();
 sky130_fd_sc_hd__nor2_4 _20614_ (.A(net318),
    .B(_08283_),
    .Y(_08294_));
 sky130_fd_sc_hd__nor2_1 _20615_ (.A(_08266_),
    .B(_08294_),
    .Y(_08295_));
 sky130_fd_sc_hd__o221ai_2 _20616_ (.A1(_12918_),
    .A2(_08284_),
    .B1(_08289_),
    .B2(_12916_),
    .C1(_08295_),
    .Y(_08296_));
 sky130_fd_sc_hd__xnor2_4 _20617_ (.A(\count_hash1[4] ),
    .B(_10351_),
    .Y(_08297_));
 sky130_fd_sc_hd__nand2_4 _20618_ (.A(_08297_),
    .B(_08266_),
    .Y(_08298_));
 sky130_fd_sc_hd__nor2_4 _20619_ (.A(net319),
    .B(_08298_),
    .Y(_08299_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_964 ();
 sky130_fd_sc_hd__nand2_2 _20621_ (.A(net319),
    .B(net290),
    .Y(_08301_));
 sky130_fd_sc_hd__o22ai_2 _20622_ (.A1(_08297_),
    .A2(_08301_),
    .B1(_08298_),
    .B2(net319),
    .Y(_08302_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_963 ();
 sky130_fd_sc_hd__nand2_8 _20624_ (.A(net318),
    .B(net319),
    .Y(_08304_));
 sky130_fd_sc_hd__nand2_1 _20625_ (.A(_12912_),
    .B(net290),
    .Y(_08305_));
 sky130_fd_sc_hd__nor2_2 _20626_ (.A(_08304_),
    .B(_08305_),
    .Y(_08306_));
 sky130_fd_sc_hd__a221oi_4 _20627_ (.A1(_12916_),
    .A2(_08299_),
    .B1(_08302_),
    .B2(_12918_),
    .C1(_08306_),
    .Y(_08307_));
 sky130_fd_sc_hd__nand2_2 _20628_ (.A(net316),
    .B(_08266_),
    .Y(_08308_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_962 ();
 sky130_fd_sc_hd__nor2_4 _20630_ (.A(_12911_),
    .B(_12916_),
    .Y(_08310_));
 sky130_fd_sc_hd__nor3_1 _20631_ (.A(net319),
    .B(_08308_),
    .C(_08310_),
    .Y(_08311_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_961 ();
 sky130_fd_sc_hd__nor2_4 _20633_ (.A(net318),
    .B(_10373_),
    .Y(_08313_));
 sky130_fd_sc_hd__nand2_1 _20634_ (.A(_12916_),
    .B(_08313_),
    .Y(_08314_));
 sky130_fd_sc_hd__nand2_4 _20635_ (.A(net318),
    .B(net290),
    .Y(_08315_));
 sky130_fd_sc_hd__nand2_1 _20636_ (.A(_12912_),
    .B(_08315_),
    .Y(_08316_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_960 ();
 sky130_fd_sc_hd__a21oi_1 _20638_ (.A1(_08314_),
    .A2(_08316_),
    .B1(_08283_),
    .Y(_08318_));
 sky130_fd_sc_hd__nor2_1 _20639_ (.A(_08311_),
    .B(_08318_),
    .Y(_08319_));
 sky130_fd_sc_hd__or2_4 _20640_ (.A(\count_hash1[6] ),
    .B(_09874_),
    .X(_08320_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_959 ();
 sky130_fd_sc_hd__nor2_4 _20642_ (.A(net349),
    .B(_08320_),
    .Y(_08322_));
 sky130_fd_sc_hd__nor2_4 _20643_ (.A(_12911_),
    .B(_12918_),
    .Y(_08323_));
 sky130_fd_sc_hd__or3_1 _20644_ (.A(_12911_),
    .B(_12912_),
    .C(_12916_),
    .X(_08324_));
 sky130_fd_sc_hd__nor2_4 _20645_ (.A(net320),
    .B(net290),
    .Y(_08325_));
 sky130_fd_sc_hd__nand2_1 _20646_ (.A(_08324_),
    .B(_08325_),
    .Y(_08326_));
 sky130_fd_sc_hd__o21ai_2 _20647_ (.A1(_08283_),
    .A2(_08323_),
    .B1(_08326_),
    .Y(_08327_));
 sky130_fd_sc_hd__nand2_8 _20648_ (.A(net318),
    .B(_08327_),
    .Y(_08328_));
 sky130_fd_sc_hd__nor2_1 _20649_ (.A(_12911_),
    .B(_12912_),
    .Y(_08329_));
 sky130_fd_sc_hd__nor2_4 _20650_ (.A(_12916_),
    .B(_12918_),
    .Y(_08330_));
 sky130_fd_sc_hd__nand2_2 _20651_ (.A(_08329_),
    .B(_08330_),
    .Y(_08331_));
 sky130_fd_sc_hd__nor2_4 _20652_ (.A(_08297_),
    .B(_10373_),
    .Y(_08332_));
 sky130_fd_sc_hd__nor2_4 _20653_ (.A(_12912_),
    .B(_12916_),
    .Y(_08333_));
 sky130_fd_sc_hd__a21oi_2 _20654_ (.A1(net320),
    .A2(_08333_),
    .B1(_08325_),
    .Y(_08334_));
 sky130_fd_sc_hd__o22ai_4 _20655_ (.A1(_08331_),
    .A2(_08332_),
    .B1(_08334_),
    .B2(_08297_),
    .Y(_08335_));
 sky130_fd_sc_hd__nand2_8 _20656_ (.A(_08328_),
    .B(_08335_),
    .Y(_08336_));
 sky130_fd_sc_hd__nand2_8 _20657_ (.A(_08322_),
    .B(_08336_),
    .Y(_08337_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_958 ();
 sky130_fd_sc_hd__a31oi_1 _20659_ (.A1(_08296_),
    .A2(_08307_),
    .A3(_08319_),
    .B1(_08337_),
    .Y(_00969_));
 sky130_fd_sc_hd__nand2_2 _20660_ (.A(_08297_),
    .B(net319),
    .Y(_08339_));
 sky130_fd_sc_hd__nand2_4 _20661_ (.A(_12911_),
    .B(_08266_),
    .Y(_08340_));
 sky130_fd_sc_hd__o21ai_2 _20662_ (.A1(_08339_),
    .A2(_08340_),
    .B1(_08336_),
    .Y(_08341_));
 sky130_fd_sc_hd__a21oi_1 _20663_ (.A1(_12916_),
    .A2(_10373_),
    .B1(_08339_),
    .Y(_08342_));
 sky130_fd_sc_hd__nor2_4 _20664_ (.A(_08297_),
    .B(_08266_),
    .Y(_08343_));
 sky130_fd_sc_hd__a21oi_1 _20665_ (.A1(net319),
    .A2(_08343_),
    .B1(_08310_),
    .Y(_08344_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_957 ();
 sky130_fd_sc_hd__a21oi_1 _20667_ (.A1(_12916_),
    .A2(_08297_),
    .B1(_12911_),
    .Y(_08346_));
 sky130_fd_sc_hd__o21ai_0 _20668_ (.A1(_08332_),
    .A2(_08346_),
    .B1(_08283_),
    .Y(_08347_));
 sky130_fd_sc_hd__o21ai_0 _20669_ (.A1(_12912_),
    .A2(_08344_),
    .B1(_08347_),
    .Y(_08348_));
 sky130_fd_sc_hd__nor2_1 _20670_ (.A(_08342_),
    .B(_08348_),
    .Y(_08349_));
 sky130_fd_sc_hd__nor2_4 _20671_ (.A(\count_hash1[6] ),
    .B(_09874_),
    .Y(_08350_));
 sky130_fd_sc_hd__o21ai_0 _20672_ (.A1(_08341_),
    .A2(_08349_),
    .B1(_08350_),
    .Y(_08351_));
 sky130_fd_sc_hd__nand2b_1 _20673_ (.A_N(net348),
    .B(_08351_),
    .Y(_00970_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_956 ();
 sky130_fd_sc_hd__and2_4 _20675_ (.A(_12918_),
    .B(net320),
    .X(_08353_));
 sky130_fd_sc_hd__a21oi_1 _20676_ (.A1(_12912_),
    .A2(_08283_),
    .B1(_08353_),
    .Y(_08354_));
 sky130_fd_sc_hd__nor2_2 _20677_ (.A(_08297_),
    .B(net319),
    .Y(_08355_));
 sky130_fd_sc_hd__nor2_4 _20678_ (.A(_08283_),
    .B(_08266_),
    .Y(_08356_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_955 ();
 sky130_fd_sc_hd__o21ai_0 _20680_ (.A1(_08355_),
    .A2(_08356_),
    .B1(_12911_),
    .Y(_08358_));
 sky130_fd_sc_hd__nor2_4 _20681_ (.A(net316),
    .B(net319),
    .Y(_08359_));
 sky130_fd_sc_hd__nor2_4 _20682_ (.A(_08297_),
    .B(_08283_),
    .Y(_08360_));
 sky130_fd_sc_hd__nor2_4 _20683_ (.A(_08359_),
    .B(_08360_),
    .Y(_08361_));
 sky130_fd_sc_hd__nand2_4 _20684_ (.A(_08297_),
    .B(net289),
    .Y(_08362_));
 sky130_fd_sc_hd__a21oi_1 _20685_ (.A1(_08283_),
    .A2(_08362_),
    .B1(_12916_),
    .Y(_08363_));
 sky130_fd_sc_hd__a21oi_1 _20686_ (.A1(_08324_),
    .A2(_08284_),
    .B1(_12918_),
    .Y(_08364_));
 sky130_fd_sc_hd__a211o_1 _20687_ (.A1(_08266_),
    .A2(_08361_),
    .B1(_08363_),
    .C1(_08364_),
    .X(_08365_));
 sky130_fd_sc_hd__nor2_4 _20688_ (.A(_08283_),
    .B(net290),
    .Y(_08366_));
 sky130_fd_sc_hd__nor2_4 _20689_ (.A(net319),
    .B(_08266_),
    .Y(_08367_));
 sky130_fd_sc_hd__a22oi_1 _20690_ (.A1(_12916_),
    .A2(_08366_),
    .B1(_08367_),
    .B2(_12912_),
    .Y(_08368_));
 sky130_fd_sc_hd__nor2_2 _20691_ (.A(net316),
    .B(_08368_),
    .Y(_08369_));
 sky130_fd_sc_hd__and2_4 _20692_ (.A(_08328_),
    .B(_08335_),
    .X(_08370_));
 sky130_fd_sc_hd__a211oi_2 _20693_ (.A1(_08332_),
    .A2(_08353_),
    .B1(_08369_),
    .C1(_08370_),
    .Y(_08371_));
 sky130_fd_sc_hd__o2111ai_1 _20694_ (.A1(_08315_),
    .A2(_08354_),
    .B1(_08358_),
    .C1(_08365_),
    .D1(_08371_),
    .Y(_08372_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_954 ();
 sky130_fd_sc_hd__a21o_1 _20696_ (.A1(_08350_),
    .A2(_08372_),
    .B1(net348),
    .X(_00971_));
 sky130_fd_sc_hd__nor2_4 _20697_ (.A(_08366_),
    .B(_08367_),
    .Y(_08374_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_953 ();
 sky130_fd_sc_hd__o22ai_1 _20699_ (.A1(_08283_),
    .A2(_08362_),
    .B1(_08374_),
    .B2(_08297_),
    .Y(_08376_));
 sky130_fd_sc_hd__nand2_4 _20700_ (.A(net319),
    .B(_08266_),
    .Y(_08377_));
 sky130_fd_sc_hd__nand2_4 _20701_ (.A(_12918_),
    .B(_08297_),
    .Y(_08378_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_952 ();
 sky130_fd_sc_hd__o22ai_1 _20703_ (.A1(net290),
    .A2(_08284_),
    .B1(_08362_),
    .B2(_08283_),
    .Y(_08380_));
 sky130_fd_sc_hd__nand2_1 _20704_ (.A(_12911_),
    .B(_08380_),
    .Y(_08381_));
 sky130_fd_sc_hd__o21ai_0 _20705_ (.A1(_08377_),
    .A2(_08378_),
    .B1(_08381_),
    .Y(_08382_));
 sky130_fd_sc_hd__a21oi_1 _20706_ (.A1(_12916_),
    .A2(_08376_),
    .B1(_08382_),
    .Y(_08383_));
 sky130_fd_sc_hd__a21oi_1 _20707_ (.A1(_12911_),
    .A2(_08359_),
    .B1(_08306_),
    .Y(_08384_));
 sky130_fd_sc_hd__a21oi_1 _20708_ (.A1(_08383_),
    .A2(_08384_),
    .B1(_08337_),
    .Y(_00972_));
 sky130_fd_sc_hd__o21ai_0 _20709_ (.A1(_08299_),
    .A2(_08360_),
    .B1(_12918_),
    .Y(_08385_));
 sky130_fd_sc_hd__o21ai_0 _20710_ (.A1(_08356_),
    .A2(_08313_),
    .B1(_12912_),
    .Y(_08386_));
 sky130_fd_sc_hd__nor2_1 _20711_ (.A(net318),
    .B(_08266_),
    .Y(_08387_));
 sky130_fd_sc_hd__o21ai_0 _20712_ (.A1(_08355_),
    .A2(_08387_),
    .B1(_12911_),
    .Y(_08388_));
 sky130_fd_sc_hd__nor2_1 _20713_ (.A(_08266_),
    .B(_08359_),
    .Y(_08389_));
 sky130_fd_sc_hd__o21ai_0 _20714_ (.A1(_08299_),
    .A2(_08389_),
    .B1(_12916_),
    .Y(_08390_));
 sky130_fd_sc_hd__nand4_1 _20715_ (.A(_08385_),
    .B(_08386_),
    .C(_08388_),
    .D(_08390_),
    .Y(_08391_));
 sky130_fd_sc_hd__o21ai_0 _20716_ (.A1(_08341_),
    .A2(_08391_),
    .B1(_08350_),
    .Y(_08392_));
 sky130_fd_sc_hd__nand2b_1 _20717_ (.A_N(net348),
    .B(_08392_),
    .Y(_00973_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_951 ();
 sky130_fd_sc_hd__nand2_2 _20719_ (.A(_08283_),
    .B(net290),
    .Y(_08394_));
 sky130_fd_sc_hd__o21ai_0 _20720_ (.A1(_08283_),
    .A2(_08298_),
    .B1(_08394_),
    .Y(_08395_));
 sky130_fd_sc_hd__a22o_1 _20721_ (.A1(_12918_),
    .A2(_08356_),
    .B1(_08374_),
    .B2(_12916_),
    .X(_08396_));
 sky130_fd_sc_hd__nand2_1 _20722_ (.A(_12911_),
    .B(net290),
    .Y(_08397_));
 sky130_fd_sc_hd__a21oi_1 _20723_ (.A1(_08378_),
    .A2(_08397_),
    .B1(net319),
    .Y(_08398_));
 sky130_fd_sc_hd__a221oi_1 _20724_ (.A1(_12912_),
    .A2(_08395_),
    .B1(_08396_),
    .B2(net316),
    .C1(_08398_),
    .Y(_08399_));
 sky130_fd_sc_hd__a21oi_1 _20725_ (.A1(_08383_),
    .A2(_08399_),
    .B1(_08337_),
    .Y(_00974_));
 sky130_fd_sc_hd__nor2_1 _20726_ (.A(_08283_),
    .B(_08330_),
    .Y(_08400_));
 sky130_fd_sc_hd__o221ai_1 _20727_ (.A1(_12916_),
    .A2(_08304_),
    .B1(_08400_),
    .B2(_12912_),
    .C1(_08389_),
    .Y(_08401_));
 sky130_fd_sc_hd__nand2_1 _20728_ (.A(_12918_),
    .B(net290),
    .Y(_08402_));
 sky130_fd_sc_hd__nand2_1 _20729_ (.A(_08340_),
    .B(_08402_),
    .Y(_08403_));
 sky130_fd_sc_hd__o21ai_2 _20730_ (.A1(_12912_),
    .A2(_08403_),
    .B1(_08359_),
    .Y(_08404_));
 sky130_fd_sc_hd__a31oi_1 _20731_ (.A1(_08328_),
    .A2(_08401_),
    .A3(_08404_),
    .B1(_08337_),
    .Y(_00975_));
 sky130_fd_sc_hd__and2_4 _20732_ (.A(_12918_),
    .B(net290),
    .X(_08405_));
 sky130_fd_sc_hd__a21oi_1 _20733_ (.A1(_12912_),
    .A2(_08266_),
    .B1(_08405_),
    .Y(_08406_));
 sky130_fd_sc_hd__o21ai_0 _20734_ (.A1(_08297_),
    .A2(_08406_),
    .B1(_08314_),
    .Y(_08407_));
 sky130_fd_sc_hd__nand2_2 _20735_ (.A(_08283_),
    .B(_08407_),
    .Y(_08408_));
 sky130_fd_sc_hd__nor2_1 _20736_ (.A(_12912_),
    .B(_12918_),
    .Y(_08409_));
 sky130_fd_sc_hd__a21oi_1 _20737_ (.A1(_08297_),
    .A2(_08409_),
    .B1(_08283_),
    .Y(_08410_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_950 ();
 sky130_fd_sc_hd__nor2_1 _20739_ (.A(_12918_),
    .B(net319),
    .Y(_08412_));
 sky130_fd_sc_hd__a21oi_1 _20740_ (.A1(net319),
    .A2(_08313_),
    .B1(_08412_),
    .Y(_08413_));
 sky130_fd_sc_hd__o21ai_0 _20741_ (.A1(_08283_),
    .A2(_08323_),
    .B1(net316),
    .Y(_08414_));
 sky130_fd_sc_hd__o221ai_1 _20742_ (.A1(_08266_),
    .A2(_08410_),
    .B1(_08413_),
    .B2(_12911_),
    .C1(_08414_),
    .Y(_08415_));
 sky130_fd_sc_hd__a21oi_2 _20743_ (.A1(_08408_),
    .A2(_08415_),
    .B1(_08337_),
    .Y(_00976_));
 sky130_fd_sc_hd__nand2_1 _20744_ (.A(net316),
    .B(_08377_),
    .Y(_08416_));
 sky130_fd_sc_hd__o21ai_0 _20745_ (.A1(_08283_),
    .A2(_08298_),
    .B1(_08416_),
    .Y(_08417_));
 sky130_fd_sc_hd__nand2_1 _20746_ (.A(_08315_),
    .B(_08298_),
    .Y(_08418_));
 sky130_fd_sc_hd__nor3_1 _20747_ (.A(_08266_),
    .B(_08330_),
    .C(_08284_),
    .Y(_08419_));
 sky130_fd_sc_hd__a31oi_1 _20748_ (.A1(_12911_),
    .A2(net320),
    .A3(_08418_),
    .B1(_08419_),
    .Y(_08420_));
 sky130_fd_sc_hd__o21ai_0 _20749_ (.A1(_08332_),
    .A2(_08356_),
    .B1(_12916_),
    .Y(_08421_));
 sky130_fd_sc_hd__o21ai_0 _20750_ (.A1(net320),
    .A2(_08313_),
    .B1(_12918_),
    .Y(_08422_));
 sky130_fd_sc_hd__nand4_1 _20751_ (.A(_08336_),
    .B(_08420_),
    .C(_08421_),
    .D(_08422_),
    .Y(_08423_));
 sky130_fd_sc_hd__a21oi_1 _20752_ (.A1(_12912_),
    .A2(_08417_),
    .B1(_08423_),
    .Y(_08424_));
 sky130_fd_sc_hd__o21bai_1 _20753_ (.A1(_08320_),
    .A2(_08424_),
    .B1_N(net348),
    .Y(_00977_));
 sky130_fd_sc_hd__nor2_2 _20754_ (.A(_08343_),
    .B(_08313_),
    .Y(_08425_));
 sky130_fd_sc_hd__nand2_1 _20755_ (.A(_08323_),
    .B(_08343_),
    .Y(_08426_));
 sky130_fd_sc_hd__o21ai_0 _20756_ (.A1(_12912_),
    .A2(net290),
    .B1(_08426_),
    .Y(_08427_));
 sky130_fd_sc_hd__or2_4 _20757_ (.A(_12912_),
    .B(_12918_),
    .X(_08428_));
 sky130_fd_sc_hd__o22ai_1 _20758_ (.A1(net316),
    .A2(_08367_),
    .B1(_08428_),
    .B2(_08355_),
    .Y(_08429_));
 sky130_fd_sc_hd__a21oi_1 _20759_ (.A1(_08283_),
    .A2(_08427_),
    .B1(_08429_),
    .Y(_08430_));
 sky130_fd_sc_hd__a221oi_1 _20760_ (.A1(_12918_),
    .A2(_08294_),
    .B1(_08425_),
    .B2(_12916_),
    .C1(_08430_),
    .Y(_08431_));
 sky130_fd_sc_hd__nor2_1 _20761_ (.A(_08337_),
    .B(_08431_),
    .Y(_00978_));
 sky130_fd_sc_hd__a21oi_1 _20762_ (.A1(_12912_),
    .A2(_08297_),
    .B1(_12916_),
    .Y(_08432_));
 sky130_fd_sc_hd__nor2_1 _20763_ (.A(net319),
    .B(_08432_),
    .Y(_08433_));
 sky130_fd_sc_hd__a211oi_1 _20764_ (.A1(_12911_),
    .A2(_08339_),
    .B1(_08433_),
    .C1(_08266_),
    .Y(_08434_));
 sky130_fd_sc_hd__a221oi_1 _20765_ (.A1(_12918_),
    .A2(_08294_),
    .B1(_08361_),
    .B2(_12912_),
    .C1(net290),
    .Y(_08435_));
 sky130_fd_sc_hd__nor2_2 _20766_ (.A(_10373_),
    .B(_08333_),
    .Y(_08436_));
 sky130_fd_sc_hd__a21oi_1 _20767_ (.A1(_08328_),
    .A2(_08333_),
    .B1(_08436_),
    .Y(_08437_));
 sky130_fd_sc_hd__nand2_1 _20768_ (.A(_08266_),
    .B(_08328_),
    .Y(_08438_));
 sky130_fd_sc_hd__o21ai_0 _20769_ (.A1(_08283_),
    .A2(_08437_),
    .B1(_08438_),
    .Y(_08439_));
 sky130_fd_sc_hd__o21ai_1 _20770_ (.A1(_08283_),
    .A2(_08362_),
    .B1(_08331_),
    .Y(_08440_));
 sky130_fd_sc_hd__a21oi_2 _20771_ (.A1(net318),
    .A2(_08439_),
    .B1(_08440_),
    .Y(_08441_));
 sky130_fd_sc_hd__o211ai_1 _20772_ (.A1(_08434_),
    .A2(_08435_),
    .B1(_08307_),
    .C1(_08441_),
    .Y(_08442_));
 sky130_fd_sc_hd__a21o_1 _20773_ (.A1(_08350_),
    .A2(_08442_),
    .B1(net348),
    .X(_00979_));
 sky130_fd_sc_hd__o21ai_0 _20774_ (.A1(net290),
    .A2(_08304_),
    .B1(_08394_),
    .Y(_08443_));
 sky130_fd_sc_hd__nand2_1 _20775_ (.A(_12912_),
    .B(_08443_),
    .Y(_08444_));
 sky130_fd_sc_hd__nand2_1 _20776_ (.A(_08359_),
    .B(_08405_),
    .Y(_08445_));
 sky130_fd_sc_hd__a21oi_1 _20777_ (.A1(net319),
    .A2(_08428_),
    .B1(_12916_),
    .Y(_08446_));
 sky130_fd_sc_hd__nor2_1 _20778_ (.A(_08362_),
    .B(_08446_),
    .Y(_08447_));
 sky130_fd_sc_hd__a31oi_1 _20779_ (.A1(_12911_),
    .A2(net316),
    .A3(_08366_),
    .B1(_08447_),
    .Y(_08448_));
 sky130_fd_sc_hd__nor2_1 _20780_ (.A(_12911_),
    .B(net319),
    .Y(_08449_));
 sky130_fd_sc_hd__nor2_1 _20781_ (.A(_12918_),
    .B(_08283_),
    .Y(_08450_));
 sky130_fd_sc_hd__nor2_1 _20782_ (.A(_08449_),
    .B(_08450_),
    .Y(_08451_));
 sky130_fd_sc_hd__o211ai_1 _20783_ (.A1(_12916_),
    .A2(_08451_),
    .B1(_08304_),
    .C1(_08266_),
    .Y(_08452_));
 sky130_fd_sc_hd__a41oi_1 _20784_ (.A1(_08444_),
    .A2(_08445_),
    .A3(_08448_),
    .A4(_08452_),
    .B1(_08337_),
    .Y(_00980_));
 sky130_fd_sc_hd__nand2_1 _20785_ (.A(_12918_),
    .B(_08266_),
    .Y(_08453_));
 sky130_fd_sc_hd__nand2_1 _20786_ (.A(_12912_),
    .B(_08374_),
    .Y(_08454_));
 sky130_fd_sc_hd__nand2_1 _20787_ (.A(_12916_),
    .B(_08356_),
    .Y(_08455_));
 sky130_fd_sc_hd__nand3_1 _20788_ (.A(_08453_),
    .B(_08454_),
    .C(_08455_),
    .Y(_08456_));
 sky130_fd_sc_hd__nand2_2 _20789_ (.A(_08297_),
    .B(_08456_),
    .Y(_08457_));
 sky130_fd_sc_hd__a21oi_1 _20790_ (.A1(_08340_),
    .A2(_08402_),
    .B1(_08283_),
    .Y(_08458_));
 sky130_fd_sc_hd__o21ai_0 _20791_ (.A1(_08436_),
    .A2(_08458_),
    .B1(net316),
    .Y(_08459_));
 sky130_fd_sc_hd__a31oi_1 _20792_ (.A1(_08296_),
    .A2(_08457_),
    .A3(_08459_),
    .B1(_08337_),
    .Y(_00981_));
 sky130_fd_sc_hd__nand2_1 _20793_ (.A(_08305_),
    .B(_08453_),
    .Y(_08460_));
 sky130_fd_sc_hd__o21ai_0 _20794_ (.A1(_12916_),
    .A2(_08460_),
    .B1(_08294_),
    .Y(_08461_));
 sky130_fd_sc_hd__o31ai_2 _20795_ (.A1(net290),
    .A2(_08304_),
    .A3(_08310_),
    .B1(_08445_),
    .Y(_08462_));
 sky130_fd_sc_hd__a221oi_1 _20796_ (.A1(_12912_),
    .A2(_08299_),
    .B1(_08451_),
    .B2(_08343_),
    .C1(_08462_),
    .Y(_08463_));
 sky130_fd_sc_hd__a31oi_1 _20797_ (.A1(_08408_),
    .A2(_08461_),
    .A3(_08463_),
    .B1(_08337_),
    .Y(_00982_));
 sky130_fd_sc_hd__nand2_1 _20798_ (.A(_12916_),
    .B(_08297_),
    .Y(_08464_));
 sky130_fd_sc_hd__nor2_1 _20799_ (.A(_12912_),
    .B(_08283_),
    .Y(_08465_));
 sky130_fd_sc_hd__a221oi_1 _20800_ (.A1(_08283_),
    .A2(_08310_),
    .B1(_08464_),
    .B2(_08465_),
    .C1(net290),
    .Y(_08466_));
 sky130_fd_sc_hd__a21oi_1 _20801_ (.A1(_12911_),
    .A2(_08284_),
    .B1(_12912_),
    .Y(_08467_));
 sky130_fd_sc_hd__nor2_1 _20802_ (.A(_12911_),
    .B(_08361_),
    .Y(_08468_));
 sky130_fd_sc_hd__nor3_1 _20803_ (.A(_08266_),
    .B(_08467_),
    .C(_08468_),
    .Y(_08469_));
 sky130_fd_sc_hd__nor2_1 _20804_ (.A(_08466_),
    .B(_08469_),
    .Y(_08470_));
 sky130_fd_sc_hd__nor2_1 _20805_ (.A(_08337_),
    .B(_08470_),
    .Y(_00983_));
 sky130_fd_sc_hd__a22oi_1 _20806_ (.A1(_12918_),
    .A2(_08360_),
    .B1(_08428_),
    .B2(_08359_),
    .Y(_08471_));
 sky130_fd_sc_hd__nand2_1 _20807_ (.A(net320),
    .B(_08333_),
    .Y(_08472_));
 sky130_fd_sc_hd__o211ai_1 _20808_ (.A1(net320),
    .A2(_08331_),
    .B1(_08472_),
    .C1(_08313_),
    .Y(_08473_));
 sky130_fd_sc_hd__inv_1 _20809_ (.A(_08455_),
    .Y(_08474_));
 sky130_fd_sc_hd__nand2_1 _20810_ (.A(net290),
    .B(_08428_),
    .Y(_08475_));
 sky130_fd_sc_hd__a21oi_1 _20811_ (.A1(_08340_),
    .A2(_08475_),
    .B1(net319),
    .Y(_08476_));
 sky130_fd_sc_hd__o21ai_0 _20812_ (.A1(_08474_),
    .A2(_08476_),
    .B1(net316),
    .Y(_08477_));
 sky130_fd_sc_hd__o2111ai_1 _20813_ (.A1(_08266_),
    .A2(_08471_),
    .B1(_08473_),
    .C1(_08477_),
    .D1(_08441_),
    .Y(_08478_));
 sky130_fd_sc_hd__a21o_1 _20814_ (.A1(_08350_),
    .A2(_08478_),
    .B1(net348),
    .X(_00984_));
 sky130_fd_sc_hd__o21ai_0 _20815_ (.A1(_12911_),
    .A2(_08405_),
    .B1(_08283_),
    .Y(_08479_));
 sky130_fd_sc_hd__o21ai_0 _20816_ (.A1(_08283_),
    .A2(_08343_),
    .B1(_12916_),
    .Y(_08480_));
 sky130_fd_sc_hd__a31oi_1 _20817_ (.A1(_08444_),
    .A2(_08479_),
    .A3(_08480_),
    .B1(_08337_),
    .Y(_00985_));
 sky130_fd_sc_hd__nor2_2 _20818_ (.A(_08266_),
    .B(_08323_),
    .Y(_08481_));
 sky130_fd_sc_hd__a21oi_1 _20819_ (.A1(_12916_),
    .A2(_08266_),
    .B1(_08481_),
    .Y(_08482_));
 sky130_fd_sc_hd__a22oi_1 _20820_ (.A1(_12911_),
    .A2(_08297_),
    .B1(_08343_),
    .B2(_12918_),
    .Y(_08483_));
 sky130_fd_sc_hd__o21ai_0 _20821_ (.A1(_08332_),
    .A2(_08294_),
    .B1(_12912_),
    .Y(_08484_));
 sky130_fd_sc_hd__o221ai_1 _20822_ (.A1(_08304_),
    .A2(_08482_),
    .B1(_08483_),
    .B2(net320),
    .C1(_08484_),
    .Y(_08485_));
 sky130_fd_sc_hd__nor3_1 _20823_ (.A(_08370_),
    .B(_08369_),
    .C(_08485_),
    .Y(_08486_));
 sky130_fd_sc_hd__o21bai_2 _20824_ (.A1(_08320_),
    .A2(_08486_),
    .B1_N(net348),
    .Y(_00986_));
 sky130_fd_sc_hd__o21ai_0 _20825_ (.A1(_08297_),
    .A2(_08330_),
    .B1(_08283_),
    .Y(_08487_));
 sky130_fd_sc_hd__nand2_1 _20826_ (.A(_08378_),
    .B(_08465_),
    .Y(_08488_));
 sky130_fd_sc_hd__o21ai_0 _20827_ (.A1(net319),
    .A2(_08308_),
    .B1(_08362_),
    .Y(_08489_));
 sky130_fd_sc_hd__a32oi_2 _20828_ (.A1(net290),
    .A2(_08487_),
    .A3(_08488_),
    .B1(_08489_),
    .B2(_12911_),
    .Y(_08490_));
 sky130_fd_sc_hd__nand2_2 _20829_ (.A(_08377_),
    .B(_08394_),
    .Y(_08491_));
 sky130_fd_sc_hd__nand3_1 _20830_ (.A(_12911_),
    .B(net316),
    .C(_08491_),
    .Y(_08492_));
 sky130_fd_sc_hd__a31oi_1 _20831_ (.A1(_08473_),
    .A2(_08490_),
    .A3(_08492_),
    .B1(_08337_),
    .Y(_00987_));
 sky130_fd_sc_hd__a22oi_1 _20832_ (.A1(_12918_),
    .A2(_08332_),
    .B1(_08425_),
    .B2(_12912_),
    .Y(_08493_));
 sky130_fd_sc_hd__nor2_1 _20833_ (.A(_08283_),
    .B(_08493_),
    .Y(_08494_));
 sky130_fd_sc_hd__nand2_1 _20834_ (.A(_12911_),
    .B(_08343_),
    .Y(_08495_));
 sky130_fd_sc_hd__nand2_1 _20835_ (.A(_12916_),
    .B(_08315_),
    .Y(_08496_));
 sky130_fd_sc_hd__a21oi_1 _20836_ (.A1(_08495_),
    .A2(_08496_),
    .B1(net319),
    .Y(_08497_));
 sky130_fd_sc_hd__a211oi_1 _20837_ (.A1(_08313_),
    .A2(_08353_),
    .B1(_08494_),
    .C1(_08497_),
    .Y(_08498_));
 sky130_fd_sc_hd__a21oi_1 _20838_ (.A1(_08404_),
    .A2(_08498_),
    .B1(_08337_),
    .Y(_00988_));
 sky130_fd_sc_hd__nand2_1 _20839_ (.A(_12911_),
    .B(_08361_),
    .Y(_08499_));
 sky130_fd_sc_hd__o21ai_0 _20840_ (.A1(_08333_),
    .A2(_08284_),
    .B1(_08499_),
    .Y(_08500_));
 sky130_fd_sc_hd__nand2_1 _20841_ (.A(_08266_),
    .B(_08500_),
    .Y(_08501_));
 sky130_fd_sc_hd__a21oi_1 _20842_ (.A1(_12918_),
    .A2(_08315_),
    .B1(_12916_),
    .Y(_08502_));
 sky130_fd_sc_hd__nor2_1 _20843_ (.A(_08325_),
    .B(_08502_),
    .Y(_08503_));
 sky130_fd_sc_hd__a21oi_1 _20844_ (.A1(_08313_),
    .A2(_08450_),
    .B1(_08355_),
    .Y(_08504_));
 sky130_fd_sc_hd__o21ai_0 _20845_ (.A1(_12912_),
    .A2(_08503_),
    .B1(_08504_),
    .Y(_08505_));
 sky130_fd_sc_hd__a21oi_2 _20846_ (.A1(_08501_),
    .A2(_08505_),
    .B1(_08337_),
    .Y(_00989_));
 sky130_fd_sc_hd__nor2_1 _20847_ (.A(_12918_),
    .B(_08297_),
    .Y(_08506_));
 sky130_fd_sc_hd__a21oi_1 _20848_ (.A1(_08297_),
    .A2(_08449_),
    .B1(_08506_),
    .Y(_08507_));
 sky130_fd_sc_hd__o21ai_0 _20849_ (.A1(net316),
    .A2(_08409_),
    .B1(net319),
    .Y(_08508_));
 sky130_fd_sc_hd__o211ai_1 _20850_ (.A1(_12916_),
    .A2(_08507_),
    .B1(_08508_),
    .C1(net290),
    .Y(_08509_));
 sky130_fd_sc_hd__a21oi_1 _20851_ (.A1(_12916_),
    .A2(net316),
    .B1(_12911_),
    .Y(_08510_));
 sky130_fd_sc_hd__or3_1 _20852_ (.A(net290),
    .B(_08359_),
    .C(_08510_),
    .X(_08511_));
 sky130_fd_sc_hd__a31oi_1 _20853_ (.A1(_08307_),
    .A2(_08509_),
    .A3(_08511_),
    .B1(_08337_),
    .Y(_00990_));
 sky130_fd_sc_hd__a222oi_1 _20854_ (.A1(_12912_),
    .A2(_08301_),
    .B1(_08366_),
    .B2(_12916_),
    .C1(_08491_),
    .C2(_12911_),
    .Y(_08512_));
 sky130_fd_sc_hd__nor2_1 _20855_ (.A(_08297_),
    .B(_08512_),
    .Y(_08513_));
 sky130_fd_sc_hd__a21oi_2 _20856_ (.A1(_12916_),
    .A2(_08299_),
    .B1(_08513_),
    .Y(_08514_));
 sky130_fd_sc_hd__a31oi_2 _20857_ (.A1(_08404_),
    .A2(_08490_),
    .A3(_08514_),
    .B1(_08337_),
    .Y(_00991_));
 sky130_fd_sc_hd__o21ai_0 _20858_ (.A1(net319),
    .A2(net290),
    .B1(_12916_),
    .Y(_08515_));
 sky130_fd_sc_hd__a21oi_1 _20859_ (.A1(_08397_),
    .A2(_08515_),
    .B1(_08297_),
    .Y(_08516_));
 sky130_fd_sc_hd__a21oi_1 _20860_ (.A1(_12912_),
    .A2(_08302_),
    .B1(_08516_),
    .Y(_08517_));
 sky130_fd_sc_hd__o211ai_1 _20861_ (.A1(_08378_),
    .A2(_08491_),
    .B1(_08517_),
    .C1(_08371_),
    .Y(_08518_));
 sky130_fd_sc_hd__a21o_1 _20862_ (.A1(_08350_),
    .A2(_08518_),
    .B1(net348),
    .X(_00992_));
 sky130_fd_sc_hd__nor2_1 _20863_ (.A(_12911_),
    .B(_08266_),
    .Y(_08519_));
 sky130_fd_sc_hd__nor2_1 _20864_ (.A(net316),
    .B(_08519_),
    .Y(_08520_));
 sky130_fd_sc_hd__o22a_1 _20865_ (.A1(_12918_),
    .A2(_08298_),
    .B1(_08520_),
    .B2(_12912_),
    .X(_08521_));
 sky130_fd_sc_hd__o211ai_1 _20866_ (.A1(_12916_),
    .A2(_08521_),
    .B1(_08308_),
    .C1(net319),
    .Y(_08522_));
 sky130_fd_sc_hd__o22ai_1 _20867_ (.A1(_12911_),
    .A2(net319),
    .B1(_08377_),
    .B2(_12918_),
    .Y(_08523_));
 sky130_fd_sc_hd__a21oi_1 _20868_ (.A1(net316),
    .A2(_08523_),
    .B1(_08367_),
    .Y(_08524_));
 sky130_fd_sc_hd__o21ai_0 _20869_ (.A1(_12918_),
    .A2(_08266_),
    .B1(net316),
    .Y(_08525_));
 sky130_fd_sc_hd__nor2_1 _20870_ (.A(_12911_),
    .B(_08283_),
    .Y(_08526_));
 sky130_fd_sc_hd__nand2_1 _20871_ (.A(_08525_),
    .B(_08526_),
    .Y(_08527_));
 sky130_fd_sc_hd__o21ai_0 _20872_ (.A1(net290),
    .A2(_08412_),
    .B1(_08297_),
    .Y(_08528_));
 sky130_fd_sc_hd__o211ai_1 _20873_ (.A1(_12912_),
    .A2(_08524_),
    .B1(_08527_),
    .C1(_08528_),
    .Y(_08529_));
 sky130_fd_sc_hd__a21oi_1 _20874_ (.A1(_08522_),
    .A2(_08529_),
    .B1(_08337_),
    .Y(_00993_));
 sky130_fd_sc_hd__nand2_1 _20875_ (.A(_12916_),
    .B(_08266_),
    .Y(_08530_));
 sky130_fd_sc_hd__and2_0 _20876_ (.A(_12912_),
    .B(net290),
    .X(_08531_));
 sky130_fd_sc_hd__o21ai_0 _20877_ (.A1(_12911_),
    .A2(_08531_),
    .B1(net318),
    .Y(_08532_));
 sky130_fd_sc_hd__a21oi_1 _20878_ (.A1(_08530_),
    .A2(_08532_),
    .B1(net320),
    .Y(_08533_));
 sky130_fd_sc_hd__nor2_1 _20879_ (.A(net290),
    .B(_08323_),
    .Y(_08534_));
 sky130_fd_sc_hd__a21oi_1 _20880_ (.A1(_12916_),
    .A2(net290),
    .B1(_08534_),
    .Y(_08535_));
 sky130_fd_sc_hd__nand2_1 _20881_ (.A(_12912_),
    .B(_08299_),
    .Y(_08536_));
 sky130_fd_sc_hd__o21ai_0 _20882_ (.A1(_08304_),
    .A2(_08535_),
    .B1(_08536_),
    .Y(_08537_));
 sky130_fd_sc_hd__nor2_1 _20883_ (.A(net320),
    .B(_08329_),
    .Y(_08538_));
 sky130_fd_sc_hd__o21ai_1 _20884_ (.A1(_08400_),
    .A2(_08538_),
    .B1(_08387_),
    .Y(_08539_));
 sky130_fd_sc_hd__nor4b_1 _20885_ (.A(_08341_),
    .B(_08533_),
    .C(_08537_),
    .D_N(_08539_),
    .Y(_08540_));
 sky130_fd_sc_hd__o21bai_1 _20886_ (.A1(_08320_),
    .A2(_08540_),
    .B1_N(net348),
    .Y(_00994_));
 sky130_fd_sc_hd__nand2_1 _20887_ (.A(_08294_),
    .B(_08436_),
    .Y(_08541_));
 sky130_fd_sc_hd__nand2_2 _20888_ (.A(_08336_),
    .B(_08541_),
    .Y(_08542_));
 sky130_fd_sc_hd__nor2_1 _20889_ (.A(_08360_),
    .B(_08432_),
    .Y(_08543_));
 sky130_fd_sc_hd__nor2_1 _20890_ (.A(_12911_),
    .B(_08543_),
    .Y(_08544_));
 sky130_fd_sc_hd__nor3_1 _20891_ (.A(_12916_),
    .B(net318),
    .C(net320),
    .Y(_08545_));
 sky130_fd_sc_hd__nor3_1 _20892_ (.A(_08266_),
    .B(_08544_),
    .C(_08545_),
    .Y(_08546_));
 sky130_fd_sc_hd__o22ai_1 _20893_ (.A1(_08378_),
    .A2(_08374_),
    .B1(_08530_),
    .B2(_08297_),
    .Y(_08547_));
 sky130_fd_sc_hd__nor4_1 _20894_ (.A(_08537_),
    .B(_08542_),
    .C(_08546_),
    .D(_08547_),
    .Y(_08548_));
 sky130_fd_sc_hd__o21bai_1 _20895_ (.A1(_08320_),
    .A2(_08548_),
    .B1_N(net348),
    .Y(_00995_));
 sky130_fd_sc_hd__o21ai_1 _20896_ (.A1(_08283_),
    .A2(_08475_),
    .B1(_08515_),
    .Y(_08549_));
 sky130_fd_sc_hd__a22oi_1 _20897_ (.A1(_08360_),
    .A2(_08481_),
    .B1(_08549_),
    .B2(_08297_),
    .Y(_08550_));
 sky130_fd_sc_hd__a21oi_2 _20898_ (.A1(_08514_),
    .A2(_08550_),
    .B1(_08337_),
    .Y(_00996_));
 sky130_fd_sc_hd__o21ai_0 _20899_ (.A1(_08531_),
    .A2(_08534_),
    .B1(_08294_),
    .Y(_08551_));
 sky130_fd_sc_hd__nor2_1 _20900_ (.A(_12916_),
    .B(_08377_),
    .Y(_08552_));
 sky130_fd_sc_hd__a21oi_1 _20901_ (.A1(_12916_),
    .A2(_08301_),
    .B1(_12911_),
    .Y(_08553_));
 sky130_fd_sc_hd__or3_4 _20902_ (.A(_08297_),
    .B(_08552_),
    .C(_08553_),
    .X(_08554_));
 sky130_fd_sc_hd__a41oi_2 _20903_ (.A1(_08473_),
    .A2(_08539_),
    .A3(_08551_),
    .A4(_08554_),
    .B1(_08337_),
    .Y(_00997_));
 sky130_fd_sc_hd__a21oi_1 _20904_ (.A1(_12916_),
    .A2(net319),
    .B1(net316),
    .Y(_08555_));
 sky130_fd_sc_hd__a21oi_1 _20905_ (.A1(net319),
    .A2(_08506_),
    .B1(_08449_),
    .Y(_08556_));
 sky130_fd_sc_hd__nor2_1 _20906_ (.A(_12912_),
    .B(_08556_),
    .Y(_08557_));
 sky130_fd_sc_hd__a21oi_1 _20907_ (.A1(_12912_),
    .A2(_08284_),
    .B1(_12911_),
    .Y(_08558_));
 sky130_fd_sc_hd__nor2_1 _20908_ (.A(_08465_),
    .B(_08558_),
    .Y(_08559_));
 sky130_fd_sc_hd__o221ai_1 _20909_ (.A1(net316),
    .A2(_08325_),
    .B1(_08559_),
    .B2(_12918_),
    .C1(_08308_),
    .Y(_08560_));
 sky130_fd_sc_hd__o311ai_2 _20910_ (.A1(net290),
    .A2(_08555_),
    .A3(_08557_),
    .B1(_08448_),
    .C1(_08560_),
    .Y(_08561_));
 sky130_fd_sc_hd__o21ai_0 _20911_ (.A1(_08341_),
    .A2(_08561_),
    .B1(_08350_),
    .Y(_08562_));
 sky130_fd_sc_hd__nand2b_1 _20912_ (.A_N(net348),
    .B(_08562_),
    .Y(_00998_));
 sky130_fd_sc_hd__a21oi_1 _20913_ (.A1(_12916_),
    .A2(_08343_),
    .B1(_12911_),
    .Y(_08563_));
 sky130_fd_sc_hd__a22oi_1 _20914_ (.A1(_12912_),
    .A2(_08343_),
    .B1(_08418_),
    .B2(_12911_),
    .Y(_08564_));
 sky130_fd_sc_hd__o21ai_0 _20915_ (.A1(net320),
    .A2(_08563_),
    .B1(_08564_),
    .Y(_08565_));
 sky130_fd_sc_hd__nor4b_1 _20916_ (.A(_08462_),
    .B(_08542_),
    .C(_08565_),
    .D_N(_08457_),
    .Y(_08566_));
 sky130_fd_sc_hd__o21bai_1 _20917_ (.A1(_08320_),
    .A2(_08566_),
    .B1_N(net348),
    .Y(_00999_));
 sky130_fd_sc_hd__a22oi_1 _20918_ (.A1(_08353_),
    .A2(_08387_),
    .B1(_08425_),
    .B2(_08538_),
    .Y(_08567_));
 sky130_fd_sc_hd__nand2_1 _20919_ (.A(_12916_),
    .B(_08380_),
    .Y(_08568_));
 sky130_fd_sc_hd__nand3_1 _20920_ (.A(_08420_),
    .B(_08567_),
    .C(_08568_),
    .Y(_08569_));
 sky130_fd_sc_hd__nor3_1 _20921_ (.A(_08494_),
    .B(_08542_),
    .C(_08569_),
    .Y(_08570_));
 sky130_fd_sc_hd__o21bai_1 _20922_ (.A1(_08320_),
    .A2(_08570_),
    .B1_N(net348),
    .Y(_01000_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_948 ();
 sky130_fd_sc_hd__nor2_4 _20925_ (.A(_12902_),
    .B(_12906_),
    .Y(_08573_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_946 ();
 sky130_fd_sc_hd__nor2_4 _20928_ (.A(_12901_),
    .B(_12904_),
    .Y(_08576_));
 sky130_fd_sc_hd__nand2_8 _20929_ (.A(_08573_),
    .B(_08576_),
    .Y(_08577_));
 sky130_fd_sc_hd__nand2_8 _20930_ (.A(_08322_),
    .B(_08577_),
    .Y(_08578_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_944 ();
 sky130_fd_sc_hd__or2_4 _20933_ (.A(_12902_),
    .B(_12906_),
    .X(_08581_));
 sky130_fd_sc_hd__nor3_4 _20934_ (.A(_12901_),
    .B(_12904_),
    .C(_08581_),
    .Y(_08582_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_940 ();
 sky130_fd_sc_hd__o21ai_0 _20939_ (.A1(_12901_),
    .A2(_12906_),
    .B1(net329),
    .Y(_08587_));
 sky130_fd_sc_hd__o31ai_1 _20940_ (.A1(net329),
    .A2(net293),
    .A3(_08582_),
    .B1(_08587_),
    .Y(_08588_));
 sky130_fd_sc_hd__nor2_4 _20941_ (.A(_12901_),
    .B(_12902_),
    .Y(_08589_));
 sky130_fd_sc_hd__nor2_1 _20942_ (.A(net338),
    .B(_08589_),
    .Y(_08590_));
 sky130_fd_sc_hd__xnor2_4 _20943_ (.A(\count_hash2[3] ),
    .B(_12908_),
    .Y(_08591_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_939 ();
 sky130_fd_sc_hd__nor2_4 _20945_ (.A(_12904_),
    .B(_12906_),
    .Y(_08593_));
 sky130_fd_sc_hd__nor2_1 _20946_ (.A(_08591_),
    .B(_08593_),
    .Y(_08594_));
 sky130_fd_sc_hd__o21ai_4 _20947_ (.A1(_08590_),
    .A2(_08594_),
    .B1(_09867_),
    .Y(_08595_));
 sky130_fd_sc_hd__nand2_4 _20948_ (.A(net329),
    .B(net533),
    .Y(_08596_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_937 ();
 sky130_fd_sc_hd__xor2_4 _20951_ (.A(\count_hash2[5] ),
    .B(_09866_),
    .X(_08599_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_935 ();
 sky130_fd_sc_hd__inv_6 _20954_ (.A(_12902_),
    .Y(_08602_));
 sky130_fd_sc_hd__nand2_2 _20955_ (.A(_08602_),
    .B(_08576_),
    .Y(_08603_));
 sky130_fd_sc_hd__a21oi_1 _20956_ (.A1(_12906_),
    .A2(_08599_),
    .B1(_08603_),
    .Y(_08604_));
 sky130_fd_sc_hd__o22ai_1 _20957_ (.A1(net329),
    .A2(_08595_),
    .B1(_08596_),
    .B2(_08604_),
    .Y(_08605_));
 sky130_fd_sc_hd__a21oi_2 _20958_ (.A1(net337),
    .A2(_08588_),
    .B1(_08605_),
    .Y(_08606_));
 sky130_fd_sc_hd__o21bai_4 _20959_ (.A1(_08578_),
    .A2(_08606_),
    .B1_N(net347),
    .Y(_01001_));
 sky130_fd_sc_hd__xnor2_4 _20960_ (.A(\count_hash2[4] ),
    .B(_09856_),
    .Y(_08607_));
 sky130_fd_sc_hd__nand2_8 _20961_ (.A(_08607_),
    .B(net294),
    .Y(_08608_));
 sky130_fd_sc_hd__nor2_4 _20962_ (.A(net338),
    .B(_08608_),
    .Y(_08609_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_934 ();
 sky130_fd_sc_hd__nand2_4 _20964_ (.A(net338),
    .B(_08599_),
    .Y(_08611_));
 sky130_fd_sc_hd__nor2_1 _20965_ (.A(_08607_),
    .B(_08611_),
    .Y(_08612_));
 sky130_fd_sc_hd__o21ai_2 _20966_ (.A1(_08609_),
    .A2(_08612_),
    .B1(_12901_),
    .Y(_08613_));
 sky130_fd_sc_hd__nand2_2 _20967_ (.A(_08591_),
    .B(_08599_),
    .Y(_08614_));
 sky130_fd_sc_hd__o21ai_0 _20968_ (.A1(_08573_),
    .A2(_08614_),
    .B1(_08595_),
    .Y(_08615_));
 sky130_fd_sc_hd__a21oi_1 _20969_ (.A1(net329),
    .A2(_08615_),
    .B1(_08582_),
    .Y(_08616_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_933 ();
 sky130_fd_sc_hd__nor2_4 _20971_ (.A(net533),
    .B(_08599_),
    .Y(_08618_));
 sky130_fd_sc_hd__nor2_1 _20972_ (.A(_12906_),
    .B(_08614_),
    .Y(_08619_));
 sky130_fd_sc_hd__nor2_1 _20973_ (.A(_08618_),
    .B(_08619_),
    .Y(_08620_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_932 ();
 sky130_fd_sc_hd__nor2_1 _20975_ (.A(_12901_),
    .B(_08611_),
    .Y(_08622_));
 sky130_fd_sc_hd__a31oi_1 _20976_ (.A1(_08602_),
    .A2(_08591_),
    .A3(_09867_),
    .B1(_08622_),
    .Y(_08623_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_931 ();
 sky130_fd_sc_hd__o221ai_2 _20978_ (.A1(_12904_),
    .A2(_08620_),
    .B1(_08623_),
    .B2(_12906_),
    .C1(_08607_),
    .Y(_08625_));
 sky130_fd_sc_hd__a31oi_4 _20979_ (.A1(_08613_),
    .A2(_08616_),
    .A3(_08625_),
    .B1(_08320_),
    .Y(_08626_));
 sky130_fd_sc_hd__or2_0 _20980_ (.A(net347),
    .B(_08626_),
    .X(_01002_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_929 ();
 sky130_fd_sc_hd__nand2_2 _20983_ (.A(net533),
    .B(_08593_),
    .Y(_08629_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_928 ();
 sky130_fd_sc_hd__nor2_4 _20985_ (.A(_12902_),
    .B(_12904_),
    .Y(_08631_));
 sky130_fd_sc_hd__nand2_1 _20986_ (.A(net338),
    .B(_08631_),
    .Y(_08632_));
 sky130_fd_sc_hd__nor2_4 _20987_ (.A(net328),
    .B(_08599_),
    .Y(_08633_));
 sky130_fd_sc_hd__o211ai_1 _20988_ (.A1(_12901_),
    .A2(_08629_),
    .B1(_08632_),
    .C1(_08633_),
    .Y(_08634_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_927 ();
 sky130_fd_sc_hd__nand2_1 _20990_ (.A(_12902_),
    .B(_08607_),
    .Y(_08636_));
 sky130_fd_sc_hd__nand2_1 _20991_ (.A(_12906_),
    .B(net328),
    .Y(_08637_));
 sky130_fd_sc_hd__nand2_1 _20992_ (.A(_08636_),
    .B(_08637_),
    .Y(_08638_));
 sky130_fd_sc_hd__nor2_4 _20993_ (.A(net533),
    .B(net294),
    .Y(_08639_));
 sky130_fd_sc_hd__o21ai_0 _20994_ (.A1(_12901_),
    .A2(_08638_),
    .B1(_08639_),
    .Y(_08640_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_924 ();
 sky130_fd_sc_hd__a21oi_1 _20998_ (.A1(_12904_),
    .A2(net294),
    .B1(_12901_),
    .Y(_08644_));
 sky130_fd_sc_hd__o21ai_0 _20999_ (.A1(_08607_),
    .A2(_08644_),
    .B1(_08602_),
    .Y(_08645_));
 sky130_fd_sc_hd__nand2_1 _21000_ (.A(net533),
    .B(_08645_),
    .Y(_08646_));
 sky130_fd_sc_hd__nand2_4 _21001_ (.A(_08607_),
    .B(_08591_),
    .Y(_08647_));
 sky130_fd_sc_hd__nand2_2 _21002_ (.A(net328),
    .B(net337),
    .Y(_08648_));
 sky130_fd_sc_hd__nor2_2 _21003_ (.A(net337),
    .B(_08593_),
    .Y(_08649_));
 sky130_fd_sc_hd__a32oi_1 _21004_ (.A1(_12901_),
    .A2(_08647_),
    .A3(_08648_),
    .B1(_08649_),
    .B2(net328),
    .Y(_08650_));
 sky130_fd_sc_hd__nand2_2 _21005_ (.A(net329),
    .B(net294),
    .Y(_08651_));
 sky130_fd_sc_hd__nor2_4 _21006_ (.A(net329),
    .B(net294),
    .Y(_08652_));
 sky130_fd_sc_hd__nand2_1 _21007_ (.A(net533),
    .B(_08652_),
    .Y(_08653_));
 sky130_fd_sc_hd__o21ai_0 _21008_ (.A1(_08591_),
    .A2(_08651_),
    .B1(_08653_),
    .Y(_08654_));
 sky130_fd_sc_hd__nand2_2 _21009_ (.A(net338),
    .B(_09867_),
    .Y(_08655_));
 sky130_fd_sc_hd__nand2_4 _21010_ (.A(_12904_),
    .B(_09857_),
    .Y(_08656_));
 sky130_fd_sc_hd__o22ai_1 _21011_ (.A1(_08655_),
    .A2(_08656_),
    .B1(_08653_),
    .B2(_08573_),
    .Y(_08657_));
 sky130_fd_sc_hd__a21oi_2 _21012_ (.A1(_12901_),
    .A2(_08654_),
    .B1(_08657_),
    .Y(_08658_));
 sky130_fd_sc_hd__nand2_4 _21013_ (.A(_12906_),
    .B(net337),
    .Y(_08659_));
 sky130_fd_sc_hd__nor3_1 _21014_ (.A(_12901_),
    .B(_12904_),
    .C(_12906_),
    .Y(_08660_));
 sky130_fd_sc_hd__a21oi_1 _21015_ (.A1(net293),
    .A2(_08659_),
    .B1(_08660_),
    .Y(_08661_));
 sky130_fd_sc_hd__nor3_1 _21016_ (.A(_12902_),
    .B(_08607_),
    .C(_08661_),
    .Y(_08662_));
 sky130_fd_sc_hd__nor2_4 _21017_ (.A(net338),
    .B(net294),
    .Y(_08663_));
 sky130_fd_sc_hd__a221oi_1 _21018_ (.A1(_12904_),
    .A2(_08663_),
    .B1(_08618_),
    .B2(_12906_),
    .C1(_09857_),
    .Y(_08664_));
 sky130_fd_sc_hd__nor2_1 _21019_ (.A(_08662_),
    .B(_08664_),
    .Y(_08665_));
 sky130_fd_sc_hd__a21oi_1 _21020_ (.A1(_08577_),
    .A2(_08639_),
    .B1(_08665_),
    .Y(_08666_));
 sky130_fd_sc_hd__o211ai_1 _21021_ (.A1(_08599_),
    .A2(_08650_),
    .B1(_08658_),
    .C1(_08666_),
    .Y(_08667_));
 sky130_fd_sc_hd__a41oi_2 _21022_ (.A1(_08634_),
    .A2(_08640_),
    .A3(_08646_),
    .A4(_08667_),
    .B1(_09875_),
    .Y(_01003_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_923 ();
 sky130_fd_sc_hd__a22oi_1 _21024_ (.A1(net533),
    .A2(_08576_),
    .B1(_08618_),
    .B2(_08607_),
    .Y(_08669_));
 sky130_fd_sc_hd__nand2_4 _21025_ (.A(net329),
    .B(_08599_),
    .Y(_08670_));
 sky130_fd_sc_hd__o21ai_0 _21026_ (.A1(net337),
    .A2(_08633_),
    .B1(_12901_),
    .Y(_08671_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_922 ();
 sky130_fd_sc_hd__nor2_4 _21028_ (.A(net328),
    .B(net533),
    .Y(_08673_));
 sky130_fd_sc_hd__o21ai_0 _21029_ (.A1(_12904_),
    .A2(net293),
    .B1(_08673_),
    .Y(_08674_));
 sky130_fd_sc_hd__nand3_1 _21030_ (.A(_08670_),
    .B(_08671_),
    .C(_08674_),
    .Y(_08675_));
 sky130_fd_sc_hd__o21ai_2 _21031_ (.A1(_12902_),
    .A2(_08669_),
    .B1(_08675_),
    .Y(_08676_));
 sky130_fd_sc_hd__nor2_1 _21032_ (.A(_08578_),
    .B(_08676_),
    .Y(_01004_));
 sky130_fd_sc_hd__a21oi_2 _21033_ (.A1(_08633_),
    .A2(_08649_),
    .B1(_08582_),
    .Y(_08677_));
 sky130_fd_sc_hd__nand2_1 _21034_ (.A(_08589_),
    .B(_08656_),
    .Y(_08678_));
 sky130_fd_sc_hd__nand2_2 _21035_ (.A(_08639_),
    .B(_08678_),
    .Y(_08679_));
 sky130_fd_sc_hd__o21ai_0 _21036_ (.A1(_08602_),
    .A2(_08673_),
    .B1(_08637_),
    .Y(_08680_));
 sky130_fd_sc_hd__or3_4 _21037_ (.A(_12902_),
    .B(_12904_),
    .C(_12906_),
    .X(_08681_));
 sky130_fd_sc_hd__a22o_1 _21038_ (.A1(_12901_),
    .A2(net533),
    .B1(_08618_),
    .B2(_08681_),
    .X(_08682_));
 sky130_fd_sc_hd__a22oi_1 _21039_ (.A1(net293),
    .A2(_08680_),
    .B1(_08682_),
    .B2(_08607_),
    .Y(_08683_));
 sky130_fd_sc_hd__a31oi_2 _21040_ (.A1(_08677_),
    .A2(_08679_),
    .A3(_08683_),
    .B1(net285),
    .Y(_01005_));
 sky130_fd_sc_hd__nand3_4 _21041_ (.A(net293),
    .B(_08673_),
    .C(_08681_),
    .Y(_08684_));
 sky130_fd_sc_hd__nand2_4 _21042_ (.A(_08647_),
    .B(_08648_),
    .Y(_08685_));
 sky130_fd_sc_hd__nor2_1 _21043_ (.A(_12901_),
    .B(_08591_),
    .Y(_08686_));
 sky130_fd_sc_hd__a21oi_1 _21044_ (.A1(_12901_),
    .A2(_08647_),
    .B1(_12902_),
    .Y(_08687_));
 sky130_fd_sc_hd__a221oi_1 _21045_ (.A1(_08591_),
    .A2(_08652_),
    .B1(_08686_),
    .B2(_08670_),
    .C1(_08687_),
    .Y(_08688_));
 sky130_fd_sc_hd__o22ai_1 _21046_ (.A1(_08599_),
    .A2(_08685_),
    .B1(_08688_),
    .B2(_12906_),
    .Y(_08689_));
 sky130_fd_sc_hd__a21oi_1 _21047_ (.A1(_08684_),
    .A2(_08689_),
    .B1(_08578_),
    .Y(_08690_));
 sky130_fd_sc_hd__or2_0 _21048_ (.A(net347),
    .B(_08690_),
    .X(_01006_));
 sky130_fd_sc_hd__nand2_1 _21049_ (.A(_08591_),
    .B(_08603_),
    .Y(_08691_));
 sky130_fd_sc_hd__nand2_8 _21050_ (.A(_08607_),
    .B(_08599_),
    .Y(_08692_));
 sky130_fd_sc_hd__a21oi_1 _21051_ (.A1(_08659_),
    .A2(_08691_),
    .B1(_08692_),
    .Y(_08693_));
 sky130_fd_sc_hd__nand2_1 _21052_ (.A(_12904_),
    .B(_08599_),
    .Y(_08694_));
 sky130_fd_sc_hd__nand2_1 _21053_ (.A(_12902_),
    .B(net329),
    .Y(_08695_));
 sky130_fd_sc_hd__nor2_4 _21054_ (.A(_08607_),
    .B(_08599_),
    .Y(_08696_));
 sky130_fd_sc_hd__nor2_2 _21055_ (.A(_08652_),
    .B(_08696_),
    .Y(_08697_));
 sky130_fd_sc_hd__a221oi_1 _21056_ (.A1(_12904_),
    .A2(_08633_),
    .B1(_08697_),
    .B2(_12901_),
    .C1(net338),
    .Y(_08698_));
 sky130_fd_sc_hd__a31oi_1 _21057_ (.A1(net338),
    .A2(_08694_),
    .A3(_08695_),
    .B1(_08698_),
    .Y(_08699_));
 sky130_fd_sc_hd__nor2_1 _21058_ (.A(_08693_),
    .B(_08699_),
    .Y(_08700_));
 sky130_fd_sc_hd__nor2_1 _21059_ (.A(_08578_),
    .B(_08700_),
    .Y(_01007_));
 sky130_fd_sc_hd__nor2_2 _21060_ (.A(_08607_),
    .B(_08591_),
    .Y(_08701_));
 sky130_fd_sc_hd__a22o_1 _21061_ (.A1(_12906_),
    .A2(_08701_),
    .B1(_08685_),
    .B2(_12902_),
    .X(_08702_));
 sky130_fd_sc_hd__nand2_1 _21062_ (.A(_08599_),
    .B(_08702_),
    .Y(_08703_));
 sky130_fd_sc_hd__o22ai_1 _21063_ (.A1(_08591_),
    .A2(_08608_),
    .B1(_08614_),
    .B2(_08607_),
    .Y(_08704_));
 sky130_fd_sc_hd__nor2_2 _21064_ (.A(_08602_),
    .B(_08591_),
    .Y(_08705_));
 sky130_fd_sc_hd__nor3_1 _21065_ (.A(net293),
    .B(_08576_),
    .C(_08596_),
    .Y(_08706_));
 sky130_fd_sc_hd__a221oi_1 _21066_ (.A1(_12906_),
    .A2(_08704_),
    .B1(_08705_),
    .B2(_08633_),
    .C1(_08706_),
    .Y(_08707_));
 sky130_fd_sc_hd__a21oi_1 _21067_ (.A1(_12901_),
    .A2(_08607_),
    .B1(net533),
    .Y(_08708_));
 sky130_fd_sc_hd__nand2_1 _21068_ (.A(_08656_),
    .B(_08708_),
    .Y(_08709_));
 sky130_fd_sc_hd__a21oi_1 _21069_ (.A1(_08608_),
    .A2(_08681_),
    .B1(_12901_),
    .Y(_08710_));
 sky130_fd_sc_hd__a21oi_1 _21070_ (.A1(_12904_),
    .A2(net294),
    .B1(_08607_),
    .Y(_08711_));
 sky130_fd_sc_hd__nor3_1 _21071_ (.A(net533),
    .B(_08710_),
    .C(_08711_),
    .Y(_08712_));
 sky130_fd_sc_hd__a31oi_2 _21072_ (.A1(_12906_),
    .A2(net294),
    .A3(_08709_),
    .B1(_08712_),
    .Y(_08713_));
 sky130_fd_sc_hd__a31oi_2 _21073_ (.A1(_08703_),
    .A2(_08707_),
    .A3(_08713_),
    .B1(_08578_),
    .Y(_08714_));
 sky130_fd_sc_hd__or2_0 _21074_ (.A(net347),
    .B(_08714_),
    .X(_01008_));
 sky130_fd_sc_hd__a21oi_1 _21075_ (.A1(_12906_),
    .A2(_08608_),
    .B1(_12902_),
    .Y(_08715_));
 sky130_fd_sc_hd__nand2_2 _21076_ (.A(_12904_),
    .B(net338),
    .Y(_08716_));
 sky130_fd_sc_hd__mux2i_1 _21077_ (.A0(_12901_),
    .A1(_12906_),
    .S(_08591_),
    .Y(_08717_));
 sky130_fd_sc_hd__o22ai_1 _21078_ (.A1(_08670_),
    .A2(_08716_),
    .B1(_08717_),
    .B2(_08608_),
    .Y(_08718_));
 sky130_fd_sc_hd__nor2_1 _21079_ (.A(_08582_),
    .B(_08718_),
    .Y(_08719_));
 sky130_fd_sc_hd__a21oi_1 _21080_ (.A1(_08602_),
    .A2(net328),
    .B1(net533),
    .Y(_08720_));
 sky130_fd_sc_hd__nand2_1 _21081_ (.A(net293),
    .B(_08596_),
    .Y(_08721_));
 sky130_fd_sc_hd__o311ai_1 _21082_ (.A1(_12906_),
    .A2(net293),
    .A3(_08720_),
    .B1(_08721_),
    .C1(_12904_),
    .Y(_08722_));
 sky130_fd_sc_hd__o311ai_2 _21083_ (.A1(_08619_),
    .A2(_08673_),
    .A3(_08715_),
    .B1(_08719_),
    .C1(_08722_),
    .Y(_08723_));
 sky130_fd_sc_hd__a21o_1 _21084_ (.A1(_08350_),
    .A2(_08723_),
    .B1(net347),
    .X(_01009_));
 sky130_fd_sc_hd__nor2_1 _21085_ (.A(_12901_),
    .B(_08581_),
    .Y(_08724_));
 sky130_fd_sc_hd__o22ai_1 _21086_ (.A1(_08573_),
    .A2(_08608_),
    .B1(_08670_),
    .B2(_08724_),
    .Y(_08725_));
 sky130_fd_sc_hd__a21oi_1 _21087_ (.A1(_12906_),
    .A2(_08607_),
    .B1(_12901_),
    .Y(_08726_));
 sky130_fd_sc_hd__nor3_1 _21088_ (.A(_12904_),
    .B(_08591_),
    .C(_08692_),
    .Y(_08727_));
 sky130_fd_sc_hd__a221oi_1 _21089_ (.A1(_08591_),
    .A2(_08692_),
    .B1(_08694_),
    .B2(_08726_),
    .C1(_08727_),
    .Y(_08728_));
 sky130_fd_sc_hd__a21oi_1 _21090_ (.A1(_08591_),
    .A2(_08725_),
    .B1(_08728_),
    .Y(_08729_));
 sky130_fd_sc_hd__o21bai_1 _21091_ (.A1(_08578_),
    .A2(_08729_),
    .B1_N(net347),
    .Y(_01010_));
 sky130_fd_sc_hd__nor2_1 _21092_ (.A(_12902_),
    .B(net293),
    .Y(_08730_));
 sky130_fd_sc_hd__a211oi_2 _21093_ (.A1(net293),
    .A2(_08660_),
    .B1(_08596_),
    .C1(_08730_),
    .Y(_08731_));
 sky130_fd_sc_hd__nor2_4 _21094_ (.A(_08582_),
    .B(_08731_),
    .Y(_08732_));
 sky130_fd_sc_hd__nor2_1 _21095_ (.A(_08631_),
    .B(_08647_),
    .Y(_08733_));
 sky130_fd_sc_hd__nor2_1 _21096_ (.A(_08573_),
    .B(_08648_),
    .Y(_08734_));
 sky130_fd_sc_hd__o21ai_0 _21097_ (.A1(_08733_),
    .A2(_08734_),
    .B1(net294),
    .Y(_08735_));
 sky130_fd_sc_hd__a41oi_2 _21098_ (.A1(_08658_),
    .A2(_08679_),
    .A3(_08732_),
    .A4(_08735_),
    .B1(_09875_),
    .Y(_01011_));
 sky130_fd_sc_hd__a21oi_4 _21099_ (.A1(_08591_),
    .A2(_08581_),
    .B1(_12904_),
    .Y(_08736_));
 sky130_fd_sc_hd__o21ai_0 _21100_ (.A1(_08692_),
    .A2(_08736_),
    .B1(_08684_),
    .Y(_08737_));
 sky130_fd_sc_hd__a21oi_1 _21101_ (.A1(_08636_),
    .A2(_08656_),
    .B1(net294),
    .Y(_08738_));
 sky130_fd_sc_hd__a21oi_1 _21102_ (.A1(_12901_),
    .A2(_08608_),
    .B1(_08738_),
    .Y(_08739_));
 sky130_fd_sc_hd__o21ai_0 _21103_ (.A1(net337),
    .A2(_08576_),
    .B1(_08659_),
    .Y(_08740_));
 sky130_fd_sc_hd__a21oi_1 _21104_ (.A1(net328),
    .A2(_08740_),
    .B1(_08733_),
    .Y(_08741_));
 sky130_fd_sc_hd__o22ai_2 _21105_ (.A1(net533),
    .A2(_08739_),
    .B1(_08741_),
    .B2(_08599_),
    .Y(_08742_));
 sky130_fd_sc_hd__nor2_2 _21106_ (.A(_08737_),
    .B(_08742_),
    .Y(_08743_));
 sky130_fd_sc_hd__nor2_4 _21107_ (.A(_08578_),
    .B(_08743_),
    .Y(_01012_));
 sky130_fd_sc_hd__o21ai_0 _21108_ (.A1(net338),
    .A2(_08651_),
    .B1(_08692_),
    .Y(_08744_));
 sky130_fd_sc_hd__o21ai_0 _21109_ (.A1(net338),
    .A2(_08577_),
    .B1(_08632_),
    .Y(_08745_));
 sky130_fd_sc_hd__o21ai_0 _21110_ (.A1(_09867_),
    .A2(_08745_),
    .B1(_08595_),
    .Y(_08746_));
 sky130_fd_sc_hd__nand2_4 _21111_ (.A(_08591_),
    .B(_09867_),
    .Y(_08747_));
 sky130_fd_sc_hd__nand3_1 _21112_ (.A(_08591_),
    .B(_09867_),
    .C(_08593_),
    .Y(_08748_));
 sky130_fd_sc_hd__a21oi_1 _21113_ (.A1(_08611_),
    .A2(_08748_),
    .B1(_12901_),
    .Y(_08749_));
 sky130_fd_sc_hd__a311oi_1 _21114_ (.A1(_08747_),
    .A2(_08611_),
    .A3(_08631_),
    .B1(_08749_),
    .C1(_09857_),
    .Y(_08750_));
 sky130_fd_sc_hd__a221oi_1 _21115_ (.A1(_12906_),
    .A2(_08744_),
    .B1(_08746_),
    .B2(_09857_),
    .C1(_08750_),
    .Y(_08751_));
 sky130_fd_sc_hd__o21bai_1 _21116_ (.A1(_08578_),
    .A2(_08751_),
    .B1_N(net349),
    .Y(_01013_));
 sky130_fd_sc_hd__nand2_1 _21117_ (.A(_12906_),
    .B(_08599_),
    .Y(_08752_));
 sky130_fd_sc_hd__nand2_1 _21118_ (.A(_12902_),
    .B(net293),
    .Y(_08753_));
 sky130_fd_sc_hd__a31oi_1 _21119_ (.A1(_08576_),
    .A2(_08752_),
    .A3(_08753_),
    .B1(_08596_),
    .Y(_08754_));
 sky130_fd_sc_hd__a21oi_1 _21120_ (.A1(_08573_),
    .A2(_08694_),
    .B1(net329),
    .Y(_08755_));
 sky130_fd_sc_hd__a21oi_1 _21121_ (.A1(_12901_),
    .A2(_08685_),
    .B1(_08705_),
    .Y(_08756_));
 sky130_fd_sc_hd__nor2_1 _21122_ (.A(_08599_),
    .B(_08756_),
    .Y(_08757_));
 sky130_fd_sc_hd__nor3_1 _21123_ (.A(_08754_),
    .B(_08755_),
    .C(_08757_),
    .Y(_08758_));
 sky130_fd_sc_hd__o21bai_1 _21124_ (.A1(_08578_),
    .A2(_08758_),
    .B1_N(net347),
    .Y(_01014_));
 sky130_fd_sc_hd__nand2_1 _21125_ (.A(_08589_),
    .B(_08618_),
    .Y(_08759_));
 sky130_fd_sc_hd__o21ai_0 _21126_ (.A1(_12904_),
    .A2(net294),
    .B1(_08759_),
    .Y(_08760_));
 sky130_fd_sc_hd__a21oi_1 _21127_ (.A1(_12901_),
    .A2(net338),
    .B1(_12902_),
    .Y(_08761_));
 sky130_fd_sc_hd__nor2_1 _21128_ (.A(_08609_),
    .B(_08761_),
    .Y(_08762_));
 sky130_fd_sc_hd__a21oi_1 _21129_ (.A1(_08652_),
    .A2(_08686_),
    .B1(_08578_),
    .Y(_08763_));
 sky130_fd_sc_hd__o21ai_0 _21130_ (.A1(_12904_),
    .A2(_08762_),
    .B1(_08763_),
    .Y(_08764_));
 sky130_fd_sc_hd__a21oi_1 _21131_ (.A1(net329),
    .A2(_08760_),
    .B1(_08764_),
    .Y(_01015_));
 sky130_fd_sc_hd__nand3_1 _21132_ (.A(_12906_),
    .B(_08607_),
    .C(net533),
    .Y(_08765_));
 sky130_fd_sc_hd__nand2_4 _21133_ (.A(_08607_),
    .B(net337),
    .Y(_08766_));
 sky130_fd_sc_hd__o22ai_1 _21134_ (.A1(_12904_),
    .A2(net338),
    .B1(_08766_),
    .B2(_12906_),
    .Y(_08767_));
 sky130_fd_sc_hd__nor2_1 _21135_ (.A(_12901_),
    .B(_08599_),
    .Y(_08768_));
 sky130_fd_sc_hd__a32oi_2 _21136_ (.A1(_08608_),
    .A2(_08716_),
    .A3(_08765_),
    .B1(_08767_),
    .B2(_08768_),
    .Y(_08769_));
 sky130_fd_sc_hd__nor3_1 _21137_ (.A(_08582_),
    .B(_08706_),
    .C(_08769_),
    .Y(_08770_));
 sky130_fd_sc_hd__a21oi_1 _21138_ (.A1(_08703_),
    .A2(_08770_),
    .B1(_09875_),
    .Y(_01016_));
 sky130_fd_sc_hd__a21oi_1 _21139_ (.A1(_12904_),
    .A2(_09857_),
    .B1(_12906_),
    .Y(_08771_));
 sky130_fd_sc_hd__nand2_1 _21140_ (.A(_12904_),
    .B(_08673_),
    .Y(_08772_));
 sky130_fd_sc_hd__o221ai_1 _21141_ (.A1(_08607_),
    .A2(_08589_),
    .B1(_08771_),
    .B2(net338),
    .C1(_08772_),
    .Y(_08773_));
 sky130_fd_sc_hd__o21ai_0 _21142_ (.A1(_08591_),
    .A2(_08692_),
    .B1(_08651_),
    .Y(_08774_));
 sky130_fd_sc_hd__a22oi_1 _21143_ (.A1(_08599_),
    .A2(_08773_),
    .B1(_08774_),
    .B2(_12901_),
    .Y(_08775_));
 sky130_fd_sc_hd__o21bai_1 _21144_ (.A1(_08578_),
    .A2(_08775_),
    .B1_N(net349),
    .Y(_01017_));
 sky130_fd_sc_hd__nor2_2 _21145_ (.A(net329),
    .B(net338),
    .Y(_08776_));
 sky130_fd_sc_hd__nor2_2 _21146_ (.A(_08607_),
    .B(net293),
    .Y(_08777_));
 sky130_fd_sc_hd__nor2_1 _21147_ (.A(_08591_),
    .B(_08633_),
    .Y(_08778_));
 sky130_fd_sc_hd__nor2_1 _21148_ (.A(_12904_),
    .B(_08607_),
    .Y(_08779_));
 sky130_fd_sc_hd__o21ai_0 _21149_ (.A1(_08599_),
    .A2(_08779_),
    .B1(_08686_),
    .Y(_08780_));
 sky130_fd_sc_hd__o21ai_0 _21150_ (.A1(_12902_),
    .A2(_08778_),
    .B1(_08780_),
    .Y(_08781_));
 sky130_fd_sc_hd__o21ai_1 _21151_ (.A1(_08612_),
    .A2(_08776_),
    .B1(_12906_),
    .Y(_08782_));
 sky130_fd_sc_hd__o311ai_0 _21152_ (.A1(_08609_),
    .A2(_08777_),
    .A3(_08781_),
    .B1(_08782_),
    .C1(_08732_),
    .Y(_08783_));
 sky130_fd_sc_hd__a21oi_1 _21153_ (.A1(_12904_),
    .A2(_08776_),
    .B1(_08783_),
    .Y(_08784_));
 sky130_fd_sc_hd__nor2_1 _21154_ (.A(_09875_),
    .B(_08784_),
    .Y(_01018_));
 sky130_fd_sc_hd__nor2_1 _21155_ (.A(_08631_),
    .B(_08766_),
    .Y(_08785_));
 sky130_fd_sc_hd__a21oi_1 _21156_ (.A1(net294),
    .A2(_08649_),
    .B1(_08785_),
    .Y(_08786_));
 sky130_fd_sc_hd__o21ai_0 _21157_ (.A1(_08633_),
    .A2(_08639_),
    .B1(_12901_),
    .Y(_08787_));
 sky130_fd_sc_hd__a31oi_1 _21158_ (.A1(_08658_),
    .A2(_08786_),
    .A3(_08787_),
    .B1(_08578_),
    .Y(_01019_));
 sky130_fd_sc_hd__a22oi_1 _21159_ (.A1(_12904_),
    .A2(_08633_),
    .B1(_08697_),
    .B2(_12902_),
    .Y(_08788_));
 sky130_fd_sc_hd__o21ai_0 _21160_ (.A1(net338),
    .A2(_08670_),
    .B1(_08766_),
    .Y(_08789_));
 sky130_fd_sc_hd__a22oi_1 _21161_ (.A1(_12906_),
    .A2(_08652_),
    .B1(_08789_),
    .B2(_12901_),
    .Y(_08790_));
 sky130_fd_sc_hd__o21ai_2 _21162_ (.A1(net338),
    .A2(_08788_),
    .B1(_08790_),
    .Y(_08791_));
 sky130_fd_sc_hd__a221oi_1 _21163_ (.A1(_12906_),
    .A2(net294),
    .B1(_08663_),
    .B2(_12904_),
    .C1(_08791_),
    .Y(_08792_));
 sky130_fd_sc_hd__nor2_1 _21164_ (.A(_08578_),
    .B(_08792_),
    .Y(_01020_));
 sky130_fd_sc_hd__nand2_1 _21165_ (.A(_08651_),
    .B(_08653_),
    .Y(_08793_));
 sky130_fd_sc_hd__nand2_2 _21166_ (.A(_08747_),
    .B(_08611_),
    .Y(_08794_));
 sky130_fd_sc_hd__nand2_1 _21167_ (.A(_12906_),
    .B(_08697_),
    .Y(_08795_));
 sky130_fd_sc_hd__nand2_1 _21168_ (.A(_12901_),
    .B(_08794_),
    .Y(_08796_));
 sky130_fd_sc_hd__nor3_1 _21169_ (.A(net294),
    .B(_08631_),
    .C(_08766_),
    .Y(_08797_));
 sky130_fd_sc_hd__a31oi_1 _21170_ (.A1(_12904_),
    .A2(_08591_),
    .A3(_08696_),
    .B1(_08797_),
    .Y(_08798_));
 sky130_fd_sc_hd__o2111ai_1 _21171_ (.A1(_08656_),
    .A2(_08794_),
    .B1(_08795_),
    .C1(_08796_),
    .D1(_08798_),
    .Y(_08799_));
 sky130_fd_sc_hd__a21oi_1 _21172_ (.A1(_12902_),
    .A2(_08793_),
    .B1(_08799_),
    .Y(_08800_));
 sky130_fd_sc_hd__o21bai_1 _21173_ (.A1(_08578_),
    .A2(_08800_),
    .B1_N(net349),
    .Y(_01021_));
 sky130_fd_sc_hd__nand2_1 _21174_ (.A(_12901_),
    .B(_08652_),
    .Y(_08801_));
 sky130_fd_sc_hd__o21ai_0 _21175_ (.A1(_08652_),
    .A2(_08696_),
    .B1(_12906_),
    .Y(_08802_));
 sky130_fd_sc_hd__a21o_4 _21176_ (.A1(_08801_),
    .A2(_08802_),
    .B1(_08591_),
    .X(_08803_));
 sky130_fd_sc_hd__o21ai_0 _21177_ (.A1(_12901_),
    .A2(_08581_),
    .B1(_08663_),
    .Y(_08804_));
 sky130_fd_sc_hd__o22ai_1 _21178_ (.A1(_08589_),
    .A2(_08647_),
    .B1(_08685_),
    .B2(_08593_),
    .Y(_08805_));
 sky130_fd_sc_hd__nand2_1 _21179_ (.A(net294),
    .B(_08805_),
    .Y(_08806_));
 sky130_fd_sc_hd__a31oi_1 _21180_ (.A1(_08803_),
    .A2(_08804_),
    .A3(_08806_),
    .B1(_08578_),
    .Y(_08807_));
 sky130_fd_sc_hd__or2_0 _21181_ (.A(net349),
    .B(_08807_),
    .X(_01022_));
 sky130_fd_sc_hd__a21oi_1 _21182_ (.A1(_12901_),
    .A2(_08591_),
    .B1(_09857_),
    .Y(_08808_));
 sky130_fd_sc_hd__o21ai_0 _21183_ (.A1(_08582_),
    .A2(_08611_),
    .B1(_08808_),
    .Y(_08809_));
 sky130_fd_sc_hd__a31oi_2 _21184_ (.A1(_12906_),
    .A2(_08747_),
    .A3(_08611_),
    .B1(_08809_),
    .Y(_08810_));
 sky130_fd_sc_hd__a22oi_1 _21185_ (.A1(_12901_),
    .A2(_08663_),
    .B1(_08655_),
    .B2(_12902_),
    .Y(_08811_));
 sky130_fd_sc_hd__nand3_2 _21186_ (.A(_09857_),
    .B(_08716_),
    .C(_08811_),
    .Y(_08812_));
 sky130_fd_sc_hd__nor3b_4 _21187_ (.A(_08810_),
    .B(_08578_),
    .C_N(_08812_),
    .Y(_01023_));
 sky130_fd_sc_hd__nand2_1 _21188_ (.A(_12904_),
    .B(_08766_),
    .Y(_08813_));
 sky130_fd_sc_hd__a22oi_1 _21189_ (.A1(_12902_),
    .A2(_08776_),
    .B1(_08701_),
    .B2(_12901_),
    .Y(_08814_));
 sky130_fd_sc_hd__a21oi_1 _21190_ (.A1(_08813_),
    .A2(_08814_),
    .B1(_08599_),
    .Y(_08815_));
 sky130_fd_sc_hd__nand2_1 _21191_ (.A(_12902_),
    .B(_08639_),
    .Y(_08816_));
 sky130_fd_sc_hd__a21oi_1 _21192_ (.A1(_08796_),
    .A2(_08816_),
    .B1(_08607_),
    .Y(_08817_));
 sky130_fd_sc_hd__nor2_1 _21193_ (.A(_08815_),
    .B(_08817_),
    .Y(_08818_));
 sky130_fd_sc_hd__o2111ai_1 _21194_ (.A1(_08692_),
    .A2(_08736_),
    .B1(_08818_),
    .C1(_08707_),
    .D1(_08577_),
    .Y(_08819_));
 sky130_fd_sc_hd__a21o_1 _21195_ (.A1(_08350_),
    .A2(_08819_),
    .B1(net349),
    .X(_01024_));
 sky130_fd_sc_hd__a21oi_1 _21196_ (.A1(_12902_),
    .A2(net294),
    .B1(_12904_),
    .Y(_08820_));
 sky130_fd_sc_hd__a21oi_1 _21197_ (.A1(_12906_),
    .A2(_08663_),
    .B1(_09857_),
    .Y(_08821_));
 sky130_fd_sc_hd__o21ai_0 _21198_ (.A1(_08591_),
    .A2(_08820_),
    .B1(_08821_),
    .Y(_08822_));
 sky130_fd_sc_hd__a32oi_1 _21199_ (.A1(_12901_),
    .A2(net338),
    .A3(net294),
    .B1(_08812_),
    .B2(_08822_),
    .Y(_08823_));
 sky130_fd_sc_hd__a21oi_1 _21200_ (.A1(_08803_),
    .A2(_08823_),
    .B1(_08578_),
    .Y(_01025_));
 sky130_fd_sc_hd__a21oi_1 _21201_ (.A1(_12901_),
    .A2(net338),
    .B1(_12904_),
    .Y(_08824_));
 sky130_fd_sc_hd__nor2_1 _21202_ (.A(_08701_),
    .B(_08824_),
    .Y(_08825_));
 sky130_fd_sc_hd__o211ai_1 _21203_ (.A1(_12906_),
    .A2(_08825_),
    .B1(_08647_),
    .C1(net293),
    .Y(_08826_));
 sky130_fd_sc_hd__nor2_1 _21204_ (.A(_12906_),
    .B(_08766_),
    .Y(_08827_));
 sky130_fd_sc_hd__a21oi_1 _21205_ (.A1(_08607_),
    .A2(_08603_),
    .B1(net337),
    .Y(_08828_));
 sky130_fd_sc_hd__or4_4 _21206_ (.A(net293),
    .B(_08827_),
    .C(_08779_),
    .D(_08828_),
    .X(_08829_));
 sky130_fd_sc_hd__a31oi_4 _21207_ (.A1(_08677_),
    .A2(_08826_),
    .A3(_08829_),
    .B1(net285),
    .Y(_01026_));
 sky130_fd_sc_hd__a21oi_1 _21208_ (.A1(_12901_),
    .A2(net293),
    .B1(_12902_),
    .Y(_08830_));
 sky130_fd_sc_hd__nor2_1 _21209_ (.A(net329),
    .B(_08830_),
    .Y(_08831_));
 sky130_fd_sc_hd__a21oi_1 _21210_ (.A1(_12906_),
    .A2(_08777_),
    .B1(_08831_),
    .Y(_08832_));
 sky130_fd_sc_hd__a22oi_1 _21211_ (.A1(_12904_),
    .A2(_08777_),
    .B1(_08692_),
    .B2(_08705_),
    .Y(_08833_));
 sky130_fd_sc_hd__o211ai_1 _21212_ (.A1(net338),
    .A2(_08832_),
    .B1(_08833_),
    .C1(_08732_),
    .Y(_08834_));
 sky130_fd_sc_hd__a21o_4 _21213_ (.A1(_08350_),
    .A2(_08834_),
    .B1(net347),
    .X(_01027_));
 sky130_fd_sc_hd__a21oi_1 _21214_ (.A1(_12901_),
    .A2(net328),
    .B1(_12904_),
    .Y(_08835_));
 sky130_fd_sc_hd__nand2_1 _21215_ (.A(_12906_),
    .B(_08673_),
    .Y(_08836_));
 sky130_fd_sc_hd__o21ai_0 _21216_ (.A1(net337),
    .A2(_08835_),
    .B1(_08836_),
    .Y(_08837_));
 sky130_fd_sc_hd__a21oi_1 _21217_ (.A1(_12906_),
    .A2(_08607_),
    .B1(_12904_),
    .Y(_08838_));
 sky130_fd_sc_hd__o21ai_0 _21218_ (.A1(_08652_),
    .A2(_08838_),
    .B1(_08602_),
    .Y(_08839_));
 sky130_fd_sc_hd__a21oi_1 _21219_ (.A1(_08602_),
    .A2(_08607_),
    .B1(net337),
    .Y(_08840_));
 sky130_fd_sc_hd__o221ai_1 _21220_ (.A1(_08607_),
    .A2(_08629_),
    .B1(_08840_),
    .B2(_12901_),
    .C1(_08766_),
    .Y(_08841_));
 sky130_fd_sc_hd__nor2_1 _21221_ (.A(_08599_),
    .B(_08841_),
    .Y(_08842_));
 sky130_fd_sc_hd__a221oi_2 _21222_ (.A1(_08599_),
    .A2(_08837_),
    .B1(_08839_),
    .B2(net337),
    .C1(_08842_),
    .Y(_08843_));
 sky130_fd_sc_hd__nor2_2 _21223_ (.A(_08578_),
    .B(_08843_),
    .Y(_01028_));
 sky130_fd_sc_hd__nand2_1 _21224_ (.A(_12904_),
    .B(_08692_),
    .Y(_08844_));
 sky130_fd_sc_hd__a311o_1 _21225_ (.A1(_08602_),
    .A2(_08801_),
    .A3(_08844_),
    .B1(net338),
    .C1(_08696_),
    .X(_08845_));
 sky130_fd_sc_hd__nor2_1 _21226_ (.A(net293),
    .B(_08576_),
    .Y(_08846_));
 sky130_fd_sc_hd__a2bb2oi_1 _21227_ (.A1_N(_12906_),
    .A2_N(_08846_),
    .B1(_08777_),
    .B2(_08576_),
    .Y(_08847_));
 sky130_fd_sc_hd__o21ai_2 _21228_ (.A1(_12902_),
    .A2(_08847_),
    .B1(_08778_),
    .Y(_08848_));
 sky130_fd_sc_hd__a31oi_4 _21229_ (.A1(_08684_),
    .A2(_08845_),
    .A3(_08848_),
    .B1(_08578_),
    .Y(_01029_));
 sky130_fd_sc_hd__a21oi_1 _21230_ (.A1(_08591_),
    .A2(_09867_),
    .B1(_08593_),
    .Y(_08849_));
 sky130_fd_sc_hd__o22ai_1 _21231_ (.A1(_12904_),
    .A2(_08655_),
    .B1(_08849_),
    .B2(_12901_),
    .Y(_08850_));
 sky130_fd_sc_hd__a21oi_1 _21232_ (.A1(_08602_),
    .A2(_08850_),
    .B1(_08622_),
    .Y(_08851_));
 sky130_fd_sc_hd__nor2_1 _21233_ (.A(net294),
    .B(_08736_),
    .Y(_08852_));
 sky130_fd_sc_hd__a21oi_1 _21234_ (.A1(_12901_),
    .A2(_08747_),
    .B1(_08852_),
    .Y(_08853_));
 sky130_fd_sc_hd__a21oi_1 _21235_ (.A1(_12904_),
    .A2(_09857_),
    .B1(_12902_),
    .Y(_08854_));
 sky130_fd_sc_hd__o221ai_1 _21236_ (.A1(_08607_),
    .A2(_08853_),
    .B1(_08854_),
    .B2(_08747_),
    .C1(_08577_),
    .Y(_08855_));
 sky130_fd_sc_hd__a21oi_1 _21237_ (.A1(_08607_),
    .A2(_08851_),
    .B1(_08855_),
    .Y(_08856_));
 sky130_fd_sc_hd__o21bai_4 _21238_ (.A1(_08320_),
    .A2(_08856_),
    .B1_N(net349),
    .Y(_01030_));
 sky130_fd_sc_hd__o21ai_0 _21239_ (.A1(_08609_),
    .A2(_08639_),
    .B1(_12902_),
    .Y(_08857_));
 sky130_fd_sc_hd__nand3_1 _21240_ (.A(_12904_),
    .B(_08599_),
    .C(_08647_),
    .Y(_08858_));
 sky130_fd_sc_hd__a21oi_1 _21241_ (.A1(_08681_),
    .A2(_08858_),
    .B1(_12901_),
    .Y(_08859_));
 sky130_fd_sc_hd__a21oi_1 _21242_ (.A1(_12901_),
    .A2(_08608_),
    .B1(_08859_),
    .Y(_08860_));
 sky130_fd_sc_hd__xnor2_1 _21243_ (.A(net329),
    .B(_08794_),
    .Y(_08861_));
 sky130_fd_sc_hd__nand2_1 _21244_ (.A(_12906_),
    .B(_08861_),
    .Y(_08862_));
 sky130_fd_sc_hd__a31oi_2 _21245_ (.A1(_08857_),
    .A2(_08860_),
    .A3(_08862_),
    .B1(_09875_),
    .Y(_01031_));
 sky130_fd_sc_hd__nor2_1 _21246_ (.A(_08659_),
    .B(_08652_),
    .Y(_08863_));
 sky130_fd_sc_hd__a2111oi_0 _21247_ (.A1(_12904_),
    .A2(_08696_),
    .B1(_08791_),
    .C1(_08863_),
    .D1(_08582_),
    .Y(_08864_));
 sky130_fd_sc_hd__nor2_1 _21248_ (.A(net285),
    .B(_08864_),
    .Y(_01032_));
 sky130_fd_sc_hd__nor2_1 _21249_ (.A(net349),
    .B(_08258_),
    .Y(_01033_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_921 ();
 sky130_fd_sc_hd__nand2_8 _21251_ (.A(_09745_),
    .B(_04784_),
    .Y(_08866_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_920 ();
 sky130_fd_sc_hd__nor2_1 _21253_ (.A(_04790_),
    .B(_08866_),
    .Y(_01034_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_919 ();
 sky130_fd_sc_hd__nor2_1 _21255_ (.A(_04871_),
    .B(_08866_),
    .Y(_01035_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_918 ();
 sky130_fd_sc_hd__nor2_1 _21257_ (.A(_04883_),
    .B(_08866_),
    .Y(_01036_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_917 ();
 sky130_fd_sc_hd__nor2_1 _21259_ (.A(_04892_),
    .B(_08866_),
    .Y(_01037_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_916 ();
 sky130_fd_sc_hd__nor2_1 _21261_ (.A(_04899_),
    .B(_08866_),
    .Y(_01038_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_915 ();
 sky130_fd_sc_hd__nor2_1 _21263_ (.A(_04906_),
    .B(_08866_),
    .Y(_01039_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_914 ();
 sky130_fd_sc_hd__nor2_1 _21265_ (.A(_04913_),
    .B(_08866_),
    .Y(_01040_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_913 ();
 sky130_fd_sc_hd__nor2_1 _21267_ (.A(_04923_),
    .B(_08866_),
    .Y(_01041_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_912 ();
 sky130_fd_sc_hd__nor2_1 _21269_ (.A(_04932_),
    .B(_08866_),
    .Y(_01042_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_911 ();
 sky130_fd_sc_hd__nor2_1 _21271_ (.A(_04939_),
    .B(_08866_),
    .Y(_01043_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_909 ();
 sky130_fd_sc_hd__nor2_1 _21274_ (.A(_04951_),
    .B(_08866_),
    .Y(_01044_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_908 ();
 sky130_fd_sc_hd__nor2_1 _21276_ (.A(_04794_),
    .B(_08866_),
    .Y(_01045_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_907 ();
 sky130_fd_sc_hd__nor2_1 _21278_ (.A(_04960_),
    .B(_08866_),
    .Y(_01046_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_906 ();
 sky130_fd_sc_hd__nor2_1 _21280_ (.A(_04974_),
    .B(_08866_),
    .Y(_01047_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_905 ();
 sky130_fd_sc_hd__nor2_1 _21282_ (.A(_04984_),
    .B(_08866_),
    .Y(_01048_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_904 ();
 sky130_fd_sc_hd__nor2_1 _21284_ (.A(_04990_),
    .B(_08866_),
    .Y(_01049_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_903 ();
 sky130_fd_sc_hd__nor2_1 _21286_ (.A(net1129),
    .B(_08866_),
    .Y(_01050_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_902 ();
 sky130_fd_sc_hd__nor2_1 _21288_ (.A(_05011_),
    .B(_08866_),
    .Y(_01051_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_901 ();
 sky130_fd_sc_hd__nor2_1 _21290_ (.A(net1139),
    .B(_08866_),
    .Y(_01052_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_900 ();
 sky130_fd_sc_hd__nor2_1 _21292_ (.A(_05029_),
    .B(_08866_),
    .Y(_01053_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_898 ();
 sky130_fd_sc_hd__nor2_1 _21295_ (.A(_05035_),
    .B(_08866_),
    .Y(_01054_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_897 ();
 sky130_fd_sc_hd__nor2_1 _21297_ (.A(_05044_),
    .B(_08866_),
    .Y(_01055_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_896 ();
 sky130_fd_sc_hd__nor2_1 _21299_ (.A(_04801_),
    .B(_08866_),
    .Y(_01056_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_895 ();
 sky130_fd_sc_hd__nor2_1 _21301_ (.A(_05060_),
    .B(_08866_),
    .Y(_01057_));
 sky130_fd_sc_hd__o21bai_1 _21302_ (.A1(_05107_),
    .A2(_05109_),
    .B1_N(_13104_),
    .Y(_08893_));
 sky130_fd_sc_hd__xnor2_1 _21303_ (.A(_05103_),
    .B(_08893_),
    .Y(_08894_));
 sky130_fd_sc_hd__mux2i_4 _21304_ (.A0(\w[62][31] ),
    .A1(_08894_),
    .S(_04797_),
    .Y(_08895_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_894 ();
 sky130_fd_sc_hd__nor2_1 _21306_ (.A(_08866_),
    .B(_08895_),
    .Y(_01058_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_893 ();
 sky130_fd_sc_hd__nor2_1 _21308_ (.A(_04808_),
    .B(_08866_),
    .Y(_01059_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_892 ();
 sky130_fd_sc_hd__nor2_1 _21310_ (.A(_04817_),
    .B(_08866_),
    .Y(_01060_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_891 ();
 sky130_fd_sc_hd__nor2_1 _21312_ (.A(_04826_),
    .B(_08866_),
    .Y(_01061_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_890 ();
 sky130_fd_sc_hd__nor2_1 _21314_ (.A(_04834_),
    .B(_08866_),
    .Y(_01062_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_889 ();
 sky130_fd_sc_hd__nor2_1 _21316_ (.A(_04843_),
    .B(_08866_),
    .Y(_01063_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_888 ();
 sky130_fd_sc_hd__nor2_1 _21318_ (.A(_04852_),
    .B(_08866_),
    .Y(_01064_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_887 ();
 sky130_fd_sc_hd__nor2_1 _21320_ (.A(_04860_),
    .B(_08866_),
    .Y(_01065_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_886 ();
 sky130_fd_sc_hd__nand2_8 _21322_ (.A(_09794_),
    .B(_05115_),
    .Y(_08905_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_885 ();
 sky130_fd_sc_hd__nor2_1 _21324_ (.A(_05118_),
    .B(_08905_),
    .Y(_01066_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_884 ();
 sky130_fd_sc_hd__nor2_1 _21326_ (.A(_05192_),
    .B(_08905_),
    .Y(_01067_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_883 ();
 sky130_fd_sc_hd__nor2_1 _21328_ (.A(_05204_),
    .B(_08905_),
    .Y(_01068_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_882 ();
 sky130_fd_sc_hd__nor2_1 _21330_ (.A(_05214_),
    .B(_08905_),
    .Y(_01069_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_881 ();
 sky130_fd_sc_hd__nor2_1 _21332_ (.A(_05221_),
    .B(_08905_),
    .Y(_01070_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_880 ();
 sky130_fd_sc_hd__nor2_1 _21334_ (.A(net1138),
    .B(_08905_),
    .Y(_01071_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_879 ();
 sky130_fd_sc_hd__nor2_1 _21336_ (.A(_05238_),
    .B(_08905_),
    .Y(_01072_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_878 ();
 sky130_fd_sc_hd__nor2_1 _21338_ (.A(_05247_),
    .B(_08905_),
    .Y(_01073_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_877 ();
 sky130_fd_sc_hd__nor2_1 _21340_ (.A(_05258_),
    .B(_08905_),
    .Y(_01074_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_876 ();
 sky130_fd_sc_hd__nor2_1 _21342_ (.A(net1136),
    .B(_08905_),
    .Y(_01075_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_874 ();
 sky130_fd_sc_hd__nor2_1 _21345_ (.A(_05280_),
    .B(_08905_),
    .Y(_01076_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_873 ();
 sky130_fd_sc_hd__nor2_1 _21347_ (.A(_05122_),
    .B(_08905_),
    .Y(_01077_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_872 ();
 sky130_fd_sc_hd__nor2_1 _21349_ (.A(_05291_),
    .B(_08905_),
    .Y(_01078_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_871 ();
 sky130_fd_sc_hd__nor2_1 _21351_ (.A(_05301_),
    .B(_08905_),
    .Y(_01079_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_870 ();
 sky130_fd_sc_hd__nor2_1 _21353_ (.A(_05309_),
    .B(_08905_),
    .Y(_01080_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_869 ();
 sky130_fd_sc_hd__nor2_1 _21355_ (.A(_05320_),
    .B(_08905_),
    .Y(_01081_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_868 ();
 sky130_fd_sc_hd__nor2_1 _21357_ (.A(net1145),
    .B(_08905_),
    .Y(_01082_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_867 ();
 sky130_fd_sc_hd__nor2_1 _21359_ (.A(_05339_),
    .B(_08905_),
    .Y(_01083_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_866 ();
 sky130_fd_sc_hd__nor2_1 _21361_ (.A(_05347_),
    .B(_08905_),
    .Y(_01084_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_865 ();
 sky130_fd_sc_hd__nor2_1 _21363_ (.A(_05358_),
    .B(_08905_),
    .Y(_01085_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_863 ();
 sky130_fd_sc_hd__nor2_1 _21366_ (.A(net1113),
    .B(_08905_),
    .Y(_01086_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_862 ();
 sky130_fd_sc_hd__nor2_1 _21368_ (.A(_05380_),
    .B(_08905_),
    .Y(_01087_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_861 ();
 sky130_fd_sc_hd__nor2_1 _21370_ (.A(_05126_),
    .B(_08905_),
    .Y(_01088_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_860 ();
 sky130_fd_sc_hd__nor2_1 _21372_ (.A(net1114),
    .B(_08905_),
    .Y(_01089_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_859 ();
 sky130_fd_sc_hd__nor2_1 _21374_ (.A(_05430_),
    .B(_08905_),
    .Y(_01090_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_858 ();
 sky130_fd_sc_hd__nor2_1 _21376_ (.A(_05132_),
    .B(_08905_),
    .Y(_01091_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_857 ();
 sky130_fd_sc_hd__nor2_1 _21378_ (.A(_05140_),
    .B(_08905_),
    .Y(_01092_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_856 ();
 sky130_fd_sc_hd__nor2_1 _21380_ (.A(_05149_),
    .B(_08905_),
    .Y(_01093_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_855 ();
 sky130_fd_sc_hd__nor2_1 _21382_ (.A(_05157_),
    .B(_08905_),
    .Y(_01094_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_854 ();
 sky130_fd_sc_hd__nor2_1 _21384_ (.A(_05166_),
    .B(_08905_),
    .Y(_01095_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_853 ();
 sky130_fd_sc_hd__nor2_1 _21386_ (.A(_05173_),
    .B(_08905_),
    .Y(_01096_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_852 ();
 sky130_fd_sc_hd__nor2_1 _21388_ (.A(_05183_),
    .B(_08905_),
    .Y(_01097_));
 sky130_fd_sc_hd__nand2_8 _21389_ (.A(_09745_),
    .B(_05433_),
    .Y(_08940_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_851 ();
 sky130_fd_sc_hd__nor2_1 _21391_ (.A(_04790_),
    .B(_08940_),
    .Y(_01098_));
 sky130_fd_sc_hd__nor2_1 _21392_ (.A(_04871_),
    .B(_08940_),
    .Y(_01099_));
 sky130_fd_sc_hd__nor2_1 _21393_ (.A(_04883_),
    .B(_08940_),
    .Y(_01100_));
 sky130_fd_sc_hd__nor2_1 _21394_ (.A(_04892_),
    .B(_08940_),
    .Y(_01101_));
 sky130_fd_sc_hd__nor2_1 _21395_ (.A(_04899_),
    .B(_08940_),
    .Y(_01102_));
 sky130_fd_sc_hd__nor2_1 _21396_ (.A(_04906_),
    .B(_08940_),
    .Y(_01103_));
 sky130_fd_sc_hd__nor2_1 _21397_ (.A(_04913_),
    .B(_08940_),
    .Y(_01104_));
 sky130_fd_sc_hd__nor2_1 _21398_ (.A(_04923_),
    .B(_08940_),
    .Y(_01105_));
 sky130_fd_sc_hd__nor2_1 _21399_ (.A(_04932_),
    .B(_08940_),
    .Y(_01106_));
 sky130_fd_sc_hd__nor2_1 _21400_ (.A(_04939_),
    .B(_08940_),
    .Y(_01107_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_850 ();
 sky130_fd_sc_hd__nor2_1 _21402_ (.A(_04951_),
    .B(_08940_),
    .Y(_01108_));
 sky130_fd_sc_hd__nor2_1 _21403_ (.A(_04794_),
    .B(_08940_),
    .Y(_01109_));
 sky130_fd_sc_hd__nor2_1 _21404_ (.A(_04960_),
    .B(_08940_),
    .Y(_01110_));
 sky130_fd_sc_hd__nor2_1 _21405_ (.A(_04974_),
    .B(_08940_),
    .Y(_01111_));
 sky130_fd_sc_hd__nor2_1 _21406_ (.A(_04984_),
    .B(_08940_),
    .Y(_01112_));
 sky130_fd_sc_hd__nor2_1 _21407_ (.A(_04990_),
    .B(_08940_),
    .Y(_01113_));
 sky130_fd_sc_hd__nor2_1 _21408_ (.A(net1129),
    .B(_08940_),
    .Y(_01114_));
 sky130_fd_sc_hd__nor2_1 _21409_ (.A(_05011_),
    .B(_08940_),
    .Y(_01115_));
 sky130_fd_sc_hd__nor2_1 _21410_ (.A(net1139),
    .B(_08940_),
    .Y(_01116_));
 sky130_fd_sc_hd__nor2_1 _21411_ (.A(_05029_),
    .B(_08940_),
    .Y(_01117_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_849 ();
 sky130_fd_sc_hd__nor2_1 _21413_ (.A(net1135),
    .B(_08940_),
    .Y(_01118_));
 sky130_fd_sc_hd__nor2_1 _21414_ (.A(_05044_),
    .B(_08940_),
    .Y(_01119_));
 sky130_fd_sc_hd__nor2_1 _21415_ (.A(_04801_),
    .B(_08940_),
    .Y(_01120_));
 sky130_fd_sc_hd__nor2_1 _21416_ (.A(_05060_),
    .B(_08940_),
    .Y(_01121_));
 sky130_fd_sc_hd__nor2_1 _21417_ (.A(_08895_),
    .B(_08940_),
    .Y(_01122_));
 sky130_fd_sc_hd__nor2_1 _21418_ (.A(_04808_),
    .B(_08940_),
    .Y(_01123_));
 sky130_fd_sc_hd__nor2_1 _21419_ (.A(_04817_),
    .B(_08940_),
    .Y(_01124_));
 sky130_fd_sc_hd__nor2_1 _21420_ (.A(_04826_),
    .B(_08940_),
    .Y(_01125_));
 sky130_fd_sc_hd__nor2_1 _21421_ (.A(_04834_),
    .B(_08940_),
    .Y(_01126_));
 sky130_fd_sc_hd__nor2_1 _21422_ (.A(_04843_),
    .B(_08940_),
    .Y(_01127_));
 sky130_fd_sc_hd__nor2_1 _21423_ (.A(_04852_),
    .B(_08940_),
    .Y(_01128_));
 sky130_fd_sc_hd__nor2_1 _21424_ (.A(_04860_),
    .B(_08940_),
    .Y(_01129_));
 sky130_fd_sc_hd__nand2_8 _21425_ (.A(_09794_),
    .B(_05474_),
    .Y(_08944_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_848 ();
 sky130_fd_sc_hd__nor2_1 _21427_ (.A(_05118_),
    .B(_08944_),
    .Y(_01130_));
 sky130_fd_sc_hd__nor2_1 _21428_ (.A(_05192_),
    .B(_08944_),
    .Y(_01131_));
 sky130_fd_sc_hd__nor2_1 _21429_ (.A(_05204_),
    .B(_08944_),
    .Y(_01132_));
 sky130_fd_sc_hd__nor2_1 _21430_ (.A(_05214_),
    .B(_08944_),
    .Y(_01133_));
 sky130_fd_sc_hd__nor2_1 _21431_ (.A(_05221_),
    .B(_08944_),
    .Y(_01134_));
 sky130_fd_sc_hd__nor2_1 _21432_ (.A(net1138),
    .B(_08944_),
    .Y(_01135_));
 sky130_fd_sc_hd__nor2_1 _21433_ (.A(_05238_),
    .B(_08944_),
    .Y(_01136_));
 sky130_fd_sc_hd__nor2_1 _21434_ (.A(net1140),
    .B(_08944_),
    .Y(_01137_));
 sky130_fd_sc_hd__nor2_1 _21435_ (.A(_05258_),
    .B(_08944_),
    .Y(_01138_));
 sky130_fd_sc_hd__nor2_1 _21436_ (.A(_05267_),
    .B(_08944_),
    .Y(_01139_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_847 ();
 sky130_fd_sc_hd__nor2_1 _21438_ (.A(_05280_),
    .B(_08944_),
    .Y(_01140_));
 sky130_fd_sc_hd__nor2_1 _21439_ (.A(_05122_),
    .B(_08944_),
    .Y(_01141_));
 sky130_fd_sc_hd__nor2_1 _21440_ (.A(_05291_),
    .B(_08944_),
    .Y(_01142_));
 sky130_fd_sc_hd__nor2_1 _21441_ (.A(_05301_),
    .B(_08944_),
    .Y(_01143_));
 sky130_fd_sc_hd__nor2_1 _21442_ (.A(_05309_),
    .B(_08944_),
    .Y(_01144_));
 sky130_fd_sc_hd__nor2_1 _21443_ (.A(_05320_),
    .B(_08944_),
    .Y(_01145_));
 sky130_fd_sc_hd__nor2_1 _21444_ (.A(net1145),
    .B(_08944_),
    .Y(_01146_));
 sky130_fd_sc_hd__nor2_1 _21445_ (.A(_05339_),
    .B(_08944_),
    .Y(_01147_));
 sky130_fd_sc_hd__nor2_1 _21446_ (.A(net1144),
    .B(_08944_),
    .Y(_01148_));
 sky130_fd_sc_hd__nor2_1 _21447_ (.A(_05358_),
    .B(_08944_),
    .Y(_01149_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_846 ();
 sky130_fd_sc_hd__nor2_1 _21449_ (.A(net1113),
    .B(_08944_),
    .Y(_01150_));
 sky130_fd_sc_hd__nor2_1 _21450_ (.A(_05380_),
    .B(_08944_),
    .Y(_01151_));
 sky130_fd_sc_hd__nor2_1 _21451_ (.A(_05126_),
    .B(_08944_),
    .Y(_01152_));
 sky130_fd_sc_hd__nor2_1 _21452_ (.A(net1114),
    .B(_08944_),
    .Y(_01153_));
 sky130_fd_sc_hd__nor2_1 _21453_ (.A(_05430_),
    .B(_08944_),
    .Y(_01154_));
 sky130_fd_sc_hd__nor2_1 _21454_ (.A(_05132_),
    .B(_08944_),
    .Y(_01155_));
 sky130_fd_sc_hd__nor2_1 _21455_ (.A(_05140_),
    .B(_08944_),
    .Y(_01156_));
 sky130_fd_sc_hd__nor2_1 _21456_ (.A(_05149_),
    .B(_08944_),
    .Y(_01157_));
 sky130_fd_sc_hd__nor2_1 _21457_ (.A(_05157_),
    .B(_08944_),
    .Y(_01158_));
 sky130_fd_sc_hd__nor2_1 _21458_ (.A(_05166_),
    .B(_08944_),
    .Y(_01159_));
 sky130_fd_sc_hd__nor2_1 _21459_ (.A(_05173_),
    .B(_08944_),
    .Y(_01160_));
 sky130_fd_sc_hd__nor2_1 _21460_ (.A(_05183_),
    .B(_08944_),
    .Y(_01161_));
 sky130_fd_sc_hd__nand2_8 _21461_ (.A(_09745_),
    .B(_05516_),
    .Y(_08948_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_845 ();
 sky130_fd_sc_hd__nor2_1 _21463_ (.A(_04790_),
    .B(_08948_),
    .Y(_01162_));
 sky130_fd_sc_hd__nor2_1 _21464_ (.A(_04871_),
    .B(_08948_),
    .Y(_01163_));
 sky130_fd_sc_hd__nor2_1 _21465_ (.A(_04883_),
    .B(_08948_),
    .Y(_01164_));
 sky130_fd_sc_hd__nor2_1 _21466_ (.A(_04892_),
    .B(_08948_),
    .Y(_01165_));
 sky130_fd_sc_hd__nor2_1 _21467_ (.A(_04899_),
    .B(_08948_),
    .Y(_01166_));
 sky130_fd_sc_hd__nor2_1 _21468_ (.A(_04906_),
    .B(_08948_),
    .Y(_01167_));
 sky130_fd_sc_hd__nor2_1 _21469_ (.A(_04913_),
    .B(_08948_),
    .Y(_01168_));
 sky130_fd_sc_hd__nor2_1 _21470_ (.A(_04923_),
    .B(_08948_),
    .Y(_01169_));
 sky130_fd_sc_hd__nor2_1 _21471_ (.A(_04932_),
    .B(_08948_),
    .Y(_01170_));
 sky130_fd_sc_hd__nor2_1 _21472_ (.A(net1142),
    .B(_08948_),
    .Y(_01171_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_844 ();
 sky130_fd_sc_hd__nor2_1 _21474_ (.A(_04951_),
    .B(_08948_),
    .Y(_01172_));
 sky130_fd_sc_hd__nor2_1 _21475_ (.A(_04794_),
    .B(_08948_),
    .Y(_01173_));
 sky130_fd_sc_hd__nor2_1 _21476_ (.A(_04960_),
    .B(_08948_),
    .Y(_01174_));
 sky130_fd_sc_hd__nor2_1 _21477_ (.A(_04974_),
    .B(_08948_),
    .Y(_01175_));
 sky130_fd_sc_hd__nor2_1 _21478_ (.A(_04984_),
    .B(_08948_),
    .Y(_01176_));
 sky130_fd_sc_hd__nor2_1 _21479_ (.A(_04990_),
    .B(_08948_),
    .Y(_01177_));
 sky130_fd_sc_hd__nor2_1 _21480_ (.A(net1128),
    .B(_08948_),
    .Y(_01178_));
 sky130_fd_sc_hd__nor2_1 _21481_ (.A(_05011_),
    .B(_08948_),
    .Y(_01179_));
 sky130_fd_sc_hd__nor2_1 _21482_ (.A(_05020_),
    .B(_08948_),
    .Y(_01180_));
 sky130_fd_sc_hd__nor2_1 _21483_ (.A(_05029_),
    .B(_08948_),
    .Y(_01181_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_843 ();
 sky130_fd_sc_hd__nor2_1 _21485_ (.A(net1135),
    .B(_08948_),
    .Y(_01182_));
 sky130_fd_sc_hd__nor2_1 _21486_ (.A(_05044_),
    .B(_08948_),
    .Y(_01183_));
 sky130_fd_sc_hd__nor2_1 _21487_ (.A(_04801_),
    .B(_08948_),
    .Y(_01184_));
 sky130_fd_sc_hd__nor2_1 _21488_ (.A(_05060_),
    .B(_08948_),
    .Y(_01185_));
 sky130_fd_sc_hd__nor2_1 _21489_ (.A(_08895_),
    .B(_08948_),
    .Y(_01186_));
 sky130_fd_sc_hd__nor2_1 _21490_ (.A(_04808_),
    .B(_08948_),
    .Y(_01187_));
 sky130_fd_sc_hd__nor2_1 _21491_ (.A(_04817_),
    .B(_08948_),
    .Y(_01188_));
 sky130_fd_sc_hd__nor2_1 _21492_ (.A(_04826_),
    .B(_08948_),
    .Y(_01189_));
 sky130_fd_sc_hd__nor2_1 _21493_ (.A(_04834_),
    .B(_08948_),
    .Y(_01190_));
 sky130_fd_sc_hd__nor2_1 _21494_ (.A(_04843_),
    .B(_08948_),
    .Y(_01191_));
 sky130_fd_sc_hd__nor2_1 _21495_ (.A(_04852_),
    .B(_08948_),
    .Y(_01192_));
 sky130_fd_sc_hd__nor2_1 _21496_ (.A(_04860_),
    .B(_08948_),
    .Y(_01193_));
 sky130_fd_sc_hd__nand2_8 _21497_ (.A(_09794_),
    .B(_05557_),
    .Y(_08952_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_842 ();
 sky130_fd_sc_hd__nor2_1 _21499_ (.A(_05118_),
    .B(_08952_),
    .Y(_01194_));
 sky130_fd_sc_hd__nor2_1 _21500_ (.A(_05192_),
    .B(_08952_),
    .Y(_01195_));
 sky130_fd_sc_hd__nor2_1 _21501_ (.A(_05204_),
    .B(_08952_),
    .Y(_01196_));
 sky130_fd_sc_hd__nor2_1 _21502_ (.A(_05214_),
    .B(_08952_),
    .Y(_01197_));
 sky130_fd_sc_hd__nor2_1 _21503_ (.A(_05221_),
    .B(_08952_),
    .Y(_01198_));
 sky130_fd_sc_hd__nor2_1 _21504_ (.A(_05228_),
    .B(_08952_),
    .Y(_01199_));
 sky130_fd_sc_hd__nor2_1 _21505_ (.A(_05238_),
    .B(_08952_),
    .Y(_01200_));
 sky130_fd_sc_hd__nor2_1 _21506_ (.A(_05247_),
    .B(_08952_),
    .Y(_01201_));
 sky130_fd_sc_hd__nor2_1 _21507_ (.A(_05258_),
    .B(_08952_),
    .Y(_01202_));
 sky130_fd_sc_hd__nor2_1 _21508_ (.A(_05267_),
    .B(_08952_),
    .Y(_01203_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_841 ();
 sky130_fd_sc_hd__nor2_1 _21510_ (.A(_05280_),
    .B(_08952_),
    .Y(_01204_));
 sky130_fd_sc_hd__nor2_1 _21511_ (.A(_05122_),
    .B(_08952_),
    .Y(_01205_));
 sky130_fd_sc_hd__nor2_1 _21512_ (.A(_05291_),
    .B(_08952_),
    .Y(_01206_));
 sky130_fd_sc_hd__nor2_1 _21513_ (.A(_05301_),
    .B(_08952_),
    .Y(_01207_));
 sky130_fd_sc_hd__nor2_1 _21514_ (.A(_05309_),
    .B(_08952_),
    .Y(_01208_));
 sky130_fd_sc_hd__nor2_1 _21515_ (.A(_05320_),
    .B(_08952_),
    .Y(_01209_));
 sky130_fd_sc_hd__nor2_1 _21516_ (.A(net1145),
    .B(_08952_),
    .Y(_01210_));
 sky130_fd_sc_hd__nor2_1 _21517_ (.A(_05339_),
    .B(_08952_),
    .Y(_01211_));
 sky130_fd_sc_hd__nor2_1 _21518_ (.A(_05347_),
    .B(_08952_),
    .Y(_01212_));
 sky130_fd_sc_hd__nor2_1 _21519_ (.A(_05358_),
    .B(_08952_),
    .Y(_01213_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_840 ();
 sky130_fd_sc_hd__nor2_1 _21521_ (.A(net1113),
    .B(_08952_),
    .Y(_01214_));
 sky130_fd_sc_hd__nor2_1 _21522_ (.A(_05380_),
    .B(_08952_),
    .Y(_01215_));
 sky130_fd_sc_hd__nor2_1 _21523_ (.A(_05126_),
    .B(_08952_),
    .Y(_01216_));
 sky130_fd_sc_hd__nor2_1 _21524_ (.A(net1114),
    .B(_08952_),
    .Y(_01217_));
 sky130_fd_sc_hd__nor2_1 _21525_ (.A(_05430_),
    .B(_08952_),
    .Y(_01218_));
 sky130_fd_sc_hd__nor2_1 _21526_ (.A(_05132_),
    .B(_08952_),
    .Y(_01219_));
 sky130_fd_sc_hd__nor2_1 _21527_ (.A(_05140_),
    .B(_08952_),
    .Y(_01220_));
 sky130_fd_sc_hd__nor2_1 _21528_ (.A(_05149_),
    .B(_08952_),
    .Y(_01221_));
 sky130_fd_sc_hd__nor2_1 _21529_ (.A(_05157_),
    .B(_08952_),
    .Y(_01222_));
 sky130_fd_sc_hd__nor2_1 _21530_ (.A(_05166_),
    .B(_08952_),
    .Y(_01223_));
 sky130_fd_sc_hd__nor2_1 _21531_ (.A(_05173_),
    .B(_08952_),
    .Y(_01224_));
 sky130_fd_sc_hd__nor2_1 _21532_ (.A(_05183_),
    .B(_08952_),
    .Y(_01225_));
 sky130_fd_sc_hd__nand2_8 _21533_ (.A(_09745_),
    .B(_05598_),
    .Y(_08956_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_839 ();
 sky130_fd_sc_hd__nor2_1 _21535_ (.A(_04790_),
    .B(_08956_),
    .Y(_01226_));
 sky130_fd_sc_hd__nor2_1 _21536_ (.A(_04871_),
    .B(_08956_),
    .Y(_01227_));
 sky130_fd_sc_hd__nor2_1 _21537_ (.A(_04883_),
    .B(_08956_),
    .Y(_01228_));
 sky130_fd_sc_hd__nor2_1 _21538_ (.A(_04892_),
    .B(_08956_),
    .Y(_01229_));
 sky130_fd_sc_hd__nor2_1 _21539_ (.A(_04899_),
    .B(_08956_),
    .Y(_01230_));
 sky130_fd_sc_hd__nor2_1 _21540_ (.A(_04906_),
    .B(_08956_),
    .Y(_01231_));
 sky130_fd_sc_hd__nor2_1 _21541_ (.A(_04913_),
    .B(_08956_),
    .Y(_01232_));
 sky130_fd_sc_hd__nor2_1 _21542_ (.A(_04923_),
    .B(_08956_),
    .Y(_01233_));
 sky130_fd_sc_hd__nor2_1 _21543_ (.A(_04932_),
    .B(_08956_),
    .Y(_01234_));
 sky130_fd_sc_hd__nor2_1 _21544_ (.A(net1142),
    .B(_08956_),
    .Y(_01235_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_838 ();
 sky130_fd_sc_hd__nor2_1 _21546_ (.A(_04951_),
    .B(_08956_),
    .Y(_01236_));
 sky130_fd_sc_hd__nor2_1 _21547_ (.A(_04794_),
    .B(_08956_),
    .Y(_01237_));
 sky130_fd_sc_hd__nor2_1 _21548_ (.A(_04960_),
    .B(_08956_),
    .Y(_01238_));
 sky130_fd_sc_hd__nor2_1 _21549_ (.A(_04974_),
    .B(_08956_),
    .Y(_01239_));
 sky130_fd_sc_hd__nor2_1 _21550_ (.A(net1137),
    .B(_08956_),
    .Y(_01240_));
 sky130_fd_sc_hd__nor2_1 _21551_ (.A(_04990_),
    .B(_08956_),
    .Y(_01241_));
 sky130_fd_sc_hd__nor2_1 _21552_ (.A(net1128),
    .B(_08956_),
    .Y(_01242_));
 sky130_fd_sc_hd__nor2_1 _21553_ (.A(_05011_),
    .B(_08956_),
    .Y(_01243_));
 sky130_fd_sc_hd__nor2_1 _21554_ (.A(net1139),
    .B(_08956_),
    .Y(_01244_));
 sky130_fd_sc_hd__nor2_1 _21555_ (.A(_05029_),
    .B(_08956_),
    .Y(_01245_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_837 ();
 sky130_fd_sc_hd__nor2_1 _21557_ (.A(_05035_),
    .B(_08956_),
    .Y(_01246_));
 sky130_fd_sc_hd__nor2_1 _21558_ (.A(_05044_),
    .B(_08956_),
    .Y(_01247_));
 sky130_fd_sc_hd__nor2_1 _21559_ (.A(_04801_),
    .B(_08956_),
    .Y(_01248_));
 sky130_fd_sc_hd__nor2_1 _21560_ (.A(_05060_),
    .B(_08956_),
    .Y(_01249_));
 sky130_fd_sc_hd__nor2_1 _21561_ (.A(_08895_),
    .B(_08956_),
    .Y(_01250_));
 sky130_fd_sc_hd__nor2_1 _21562_ (.A(_04808_),
    .B(_08956_),
    .Y(_01251_));
 sky130_fd_sc_hd__nor2_1 _21563_ (.A(_04817_),
    .B(_08956_),
    .Y(_01252_));
 sky130_fd_sc_hd__nor2_1 _21564_ (.A(_04826_),
    .B(_08956_),
    .Y(_01253_));
 sky130_fd_sc_hd__nor2_1 _21565_ (.A(_04834_),
    .B(_08956_),
    .Y(_01254_));
 sky130_fd_sc_hd__nor2_1 _21566_ (.A(_04843_),
    .B(_08956_),
    .Y(_01255_));
 sky130_fd_sc_hd__nor2_1 _21567_ (.A(_04852_),
    .B(_08956_),
    .Y(_01256_));
 sky130_fd_sc_hd__nor2_1 _21568_ (.A(_04860_),
    .B(_08956_),
    .Y(_01257_));
 sky130_fd_sc_hd__or3_4 _21569_ (.A(net1039),
    .B(_09793_),
    .C(_09803_),
    .X(_08960_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_835 ();
 sky130_fd_sc_hd__nor2_1 _21572_ (.A(_05118_),
    .B(_08960_),
    .Y(_01258_));
 sky130_fd_sc_hd__nor2_1 _21573_ (.A(_05192_),
    .B(_08960_),
    .Y(_01259_));
 sky130_fd_sc_hd__nor2_1 _21574_ (.A(_05204_),
    .B(_08960_),
    .Y(_01260_));
 sky130_fd_sc_hd__nor2_1 _21575_ (.A(_05214_),
    .B(_08960_),
    .Y(_01261_));
 sky130_fd_sc_hd__nor2_1 _21576_ (.A(_05221_),
    .B(_08960_),
    .Y(_01262_));
 sky130_fd_sc_hd__nor2_1 _21577_ (.A(_05228_),
    .B(_08960_),
    .Y(_01263_));
 sky130_fd_sc_hd__nor2_1 _21578_ (.A(_05238_),
    .B(_08960_),
    .Y(_01264_));
 sky130_fd_sc_hd__nor2_1 _21579_ (.A(_05247_),
    .B(_08960_),
    .Y(_01265_));
 sky130_fd_sc_hd__nor2_1 _21580_ (.A(_05258_),
    .B(_08960_),
    .Y(_01266_));
 sky130_fd_sc_hd__nor2_1 _21581_ (.A(net1136),
    .B(_08960_),
    .Y(_01267_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_834 ();
 sky130_fd_sc_hd__nor2_1 _21583_ (.A(_05280_),
    .B(_08960_),
    .Y(_01268_));
 sky130_fd_sc_hd__nor2_1 _21584_ (.A(_05122_),
    .B(_08960_),
    .Y(_01269_));
 sky130_fd_sc_hd__nor2_1 _21585_ (.A(_05291_),
    .B(_08960_),
    .Y(_01270_));
 sky130_fd_sc_hd__nor2_1 _21586_ (.A(_05301_),
    .B(_08960_),
    .Y(_01271_));
 sky130_fd_sc_hd__nor2_1 _21587_ (.A(_05309_),
    .B(_08960_),
    .Y(_01272_));
 sky130_fd_sc_hd__nor2_1 _21588_ (.A(_05320_),
    .B(_08960_),
    .Y(_01273_));
 sky130_fd_sc_hd__nor2_1 _21589_ (.A(net1145),
    .B(_08960_),
    .Y(_01274_));
 sky130_fd_sc_hd__nor2_1 _21590_ (.A(_05339_),
    .B(_08960_),
    .Y(_01275_));
 sky130_fd_sc_hd__nor2_1 _21591_ (.A(net1144),
    .B(_08960_),
    .Y(_01276_));
 sky130_fd_sc_hd__nor2_1 _21592_ (.A(_05358_),
    .B(_08960_),
    .Y(_01277_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_833 ();
 sky130_fd_sc_hd__nor2_1 _21594_ (.A(net1141),
    .B(_08960_),
    .Y(_01278_));
 sky130_fd_sc_hd__nor2_1 _21595_ (.A(_05380_),
    .B(_08960_),
    .Y(_01279_));
 sky130_fd_sc_hd__nor2_1 _21596_ (.A(_05126_),
    .B(_08960_),
    .Y(_01280_));
 sky130_fd_sc_hd__nor2_1 _21597_ (.A(net1143),
    .B(_08960_),
    .Y(_01281_));
 sky130_fd_sc_hd__nor2_1 _21598_ (.A(_05430_),
    .B(_08960_),
    .Y(_01282_));
 sky130_fd_sc_hd__nor2_1 _21599_ (.A(_05132_),
    .B(_08960_),
    .Y(_01283_));
 sky130_fd_sc_hd__nor2_1 _21600_ (.A(_05140_),
    .B(_08960_),
    .Y(_01284_));
 sky130_fd_sc_hd__nor2_1 _21601_ (.A(_05149_),
    .B(_08960_),
    .Y(_01285_));
 sky130_fd_sc_hd__nor2_1 _21602_ (.A(_05157_),
    .B(_08960_),
    .Y(_01286_));
 sky130_fd_sc_hd__nor2_1 _21603_ (.A(_05166_),
    .B(_08960_),
    .Y(_01287_));
 sky130_fd_sc_hd__nor2_1 _21604_ (.A(_05173_),
    .B(_08960_),
    .Y(_01288_));
 sky130_fd_sc_hd__nor2_1 _21605_ (.A(_05183_),
    .B(_08960_),
    .Y(_01289_));
 sky130_fd_sc_hd__nand2_8 _21606_ (.A(_09751_),
    .B(_04784_),
    .Y(_08965_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_832 ();
 sky130_fd_sc_hd__nor2_1 _21608_ (.A(_04790_),
    .B(_08965_),
    .Y(_01290_));
 sky130_fd_sc_hd__nor2_1 _21609_ (.A(_04871_),
    .B(_08965_),
    .Y(_01291_));
 sky130_fd_sc_hd__nor2_1 _21610_ (.A(_04883_),
    .B(_08965_),
    .Y(_01292_));
 sky130_fd_sc_hd__nor2_1 _21611_ (.A(_04892_),
    .B(_08965_),
    .Y(_01293_));
 sky130_fd_sc_hd__nor2_1 _21612_ (.A(_04899_),
    .B(_08965_),
    .Y(_01294_));
 sky130_fd_sc_hd__nor2_1 _21613_ (.A(_04906_),
    .B(_08965_),
    .Y(_01295_));
 sky130_fd_sc_hd__nor2_1 _21614_ (.A(_04913_),
    .B(_08965_),
    .Y(_01296_));
 sky130_fd_sc_hd__nor2_1 _21615_ (.A(_04923_),
    .B(_08965_),
    .Y(_01297_));
 sky130_fd_sc_hd__nor2_1 _21616_ (.A(_04932_),
    .B(_08965_),
    .Y(_01298_));
 sky130_fd_sc_hd__nor2_1 _21617_ (.A(_04939_),
    .B(_08965_),
    .Y(_01299_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_831 ();
 sky130_fd_sc_hd__nor2_1 _21619_ (.A(_04951_),
    .B(_08965_),
    .Y(_01300_));
 sky130_fd_sc_hd__nor2_1 _21620_ (.A(_04794_),
    .B(_08965_),
    .Y(_01301_));
 sky130_fd_sc_hd__nor2_1 _21621_ (.A(_04960_),
    .B(_08965_),
    .Y(_01302_));
 sky130_fd_sc_hd__nor2_1 _21622_ (.A(_04974_),
    .B(_08965_),
    .Y(_01303_));
 sky130_fd_sc_hd__nor2_1 _21623_ (.A(_04984_),
    .B(_08965_),
    .Y(_01304_));
 sky130_fd_sc_hd__nor2_1 _21624_ (.A(_04990_),
    .B(_08965_),
    .Y(_01305_));
 sky130_fd_sc_hd__nor2_1 _21625_ (.A(net1129),
    .B(_08965_),
    .Y(_01306_));
 sky130_fd_sc_hd__nor2_1 _21626_ (.A(_05011_),
    .B(_08965_),
    .Y(_01307_));
 sky130_fd_sc_hd__nor2_1 _21627_ (.A(net1139),
    .B(_08965_),
    .Y(_01308_));
 sky130_fd_sc_hd__nor2_1 _21628_ (.A(_05029_),
    .B(_08965_),
    .Y(_01309_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_830 ();
 sky130_fd_sc_hd__nor2_1 _21630_ (.A(net1135),
    .B(_08965_),
    .Y(_01310_));
 sky130_fd_sc_hd__nor2_1 _21631_ (.A(_05044_),
    .B(_08965_),
    .Y(_01311_));
 sky130_fd_sc_hd__nor2_1 _21632_ (.A(_04801_),
    .B(_08965_),
    .Y(_01312_));
 sky130_fd_sc_hd__nor2_1 _21633_ (.A(_05060_),
    .B(_08965_),
    .Y(_01313_));
 sky130_fd_sc_hd__nor2_1 _21634_ (.A(_08895_),
    .B(_08965_),
    .Y(_01314_));
 sky130_fd_sc_hd__nor2_1 _21635_ (.A(_04808_),
    .B(_08965_),
    .Y(_01315_));
 sky130_fd_sc_hd__nor2_1 _21636_ (.A(_04817_),
    .B(_08965_),
    .Y(_01316_));
 sky130_fd_sc_hd__nor2_1 _21637_ (.A(_04826_),
    .B(_08965_),
    .Y(_01317_));
 sky130_fd_sc_hd__nor2_1 _21638_ (.A(_04834_),
    .B(_08965_),
    .Y(_01318_));
 sky130_fd_sc_hd__nor2_1 _21639_ (.A(_04843_),
    .B(_08965_),
    .Y(_01319_));
 sky130_fd_sc_hd__nor2_1 _21640_ (.A(_04852_),
    .B(_08965_),
    .Y(_01320_));
 sky130_fd_sc_hd__nor2_1 _21641_ (.A(_04860_),
    .B(_08965_),
    .Y(_01321_));
 sky130_fd_sc_hd__nand2_8 _21642_ (.A(_09805_),
    .B(_05115_),
    .Y(_08969_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_829 ();
 sky130_fd_sc_hd__nor2_1 _21644_ (.A(_05118_),
    .B(_08969_),
    .Y(_01322_));
 sky130_fd_sc_hd__nor2_1 _21645_ (.A(_05192_),
    .B(_08969_),
    .Y(_01323_));
 sky130_fd_sc_hd__nor2_1 _21646_ (.A(_05204_),
    .B(_08969_),
    .Y(_01324_));
 sky130_fd_sc_hd__nor2_1 _21647_ (.A(_05214_),
    .B(_08969_),
    .Y(_01325_));
 sky130_fd_sc_hd__nor2_1 _21648_ (.A(_05221_),
    .B(_08969_),
    .Y(_01326_));
 sky130_fd_sc_hd__nor2_1 _21649_ (.A(net1138),
    .B(_08969_),
    .Y(_01327_));
 sky130_fd_sc_hd__nor2_1 _21650_ (.A(_05238_),
    .B(_08969_),
    .Y(_01328_));
 sky130_fd_sc_hd__nor2_1 _21651_ (.A(net1140),
    .B(_08969_),
    .Y(_01329_));
 sky130_fd_sc_hd__nor2_1 _21652_ (.A(_05258_),
    .B(_08969_),
    .Y(_01330_));
 sky130_fd_sc_hd__nor2_1 _21653_ (.A(net1136),
    .B(_08969_),
    .Y(_01331_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_828 ();
 sky130_fd_sc_hd__nor2_1 _21655_ (.A(_05280_),
    .B(_08969_),
    .Y(_01332_));
 sky130_fd_sc_hd__nor2_1 _21656_ (.A(_05122_),
    .B(_08969_),
    .Y(_01333_));
 sky130_fd_sc_hd__nor2_1 _21657_ (.A(_05291_),
    .B(_08969_),
    .Y(_01334_));
 sky130_fd_sc_hd__nor2_1 _21658_ (.A(_05301_),
    .B(_08969_),
    .Y(_01335_));
 sky130_fd_sc_hd__nor2_1 _21659_ (.A(_05309_),
    .B(_08969_),
    .Y(_01336_));
 sky130_fd_sc_hd__nor2_1 _21660_ (.A(_05320_),
    .B(_08969_),
    .Y(_01337_));
 sky130_fd_sc_hd__nor2_1 _21661_ (.A(net1145),
    .B(_08969_),
    .Y(_01338_));
 sky130_fd_sc_hd__nor2_1 _21662_ (.A(_05339_),
    .B(_08969_),
    .Y(_01339_));
 sky130_fd_sc_hd__nor2_1 _21663_ (.A(_05347_),
    .B(_08969_),
    .Y(_01340_));
 sky130_fd_sc_hd__nor2_1 _21664_ (.A(_05358_),
    .B(_08969_),
    .Y(_01341_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_827 ();
 sky130_fd_sc_hd__nor2_1 _21666_ (.A(net1141),
    .B(_08969_),
    .Y(_01342_));
 sky130_fd_sc_hd__nor2_1 _21667_ (.A(_05380_),
    .B(_08969_),
    .Y(_01343_));
 sky130_fd_sc_hd__nor2_1 _21668_ (.A(_05126_),
    .B(_08969_),
    .Y(_01344_));
 sky130_fd_sc_hd__nor2_1 _21669_ (.A(net1143),
    .B(_08969_),
    .Y(_01345_));
 sky130_fd_sc_hd__nor2_1 _21670_ (.A(_05430_),
    .B(_08969_),
    .Y(_01346_));
 sky130_fd_sc_hd__nor2_1 _21671_ (.A(_05132_),
    .B(_08969_),
    .Y(_01347_));
 sky130_fd_sc_hd__nor2_1 _21672_ (.A(_05140_),
    .B(_08969_),
    .Y(_01348_));
 sky130_fd_sc_hd__nor2_1 _21673_ (.A(_05149_),
    .B(_08969_),
    .Y(_01349_));
 sky130_fd_sc_hd__nor2_1 _21674_ (.A(_05157_),
    .B(_08969_),
    .Y(_01350_));
 sky130_fd_sc_hd__nor2_1 _21675_ (.A(_05166_),
    .B(_08969_),
    .Y(_01351_));
 sky130_fd_sc_hd__nor2_1 _21676_ (.A(_05173_),
    .B(_08969_),
    .Y(_01352_));
 sky130_fd_sc_hd__nor2_1 _21677_ (.A(_05183_),
    .B(_08969_),
    .Y(_01353_));
 sky130_fd_sc_hd__nand2_8 _21678_ (.A(_09751_),
    .B(_05433_),
    .Y(_08973_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_826 ();
 sky130_fd_sc_hd__nor2_1 _21680_ (.A(_04790_),
    .B(_08973_),
    .Y(_01354_));
 sky130_fd_sc_hd__nor2_1 _21681_ (.A(_04871_),
    .B(_08973_),
    .Y(_01355_));
 sky130_fd_sc_hd__nor2_1 _21682_ (.A(_04883_),
    .B(_08973_),
    .Y(_01356_));
 sky130_fd_sc_hd__nor2_1 _21683_ (.A(_04892_),
    .B(_08973_),
    .Y(_01357_));
 sky130_fd_sc_hd__nor2_1 _21684_ (.A(_04899_),
    .B(_08973_),
    .Y(_01358_));
 sky130_fd_sc_hd__nor2_1 _21685_ (.A(_04906_),
    .B(_08973_),
    .Y(_01359_));
 sky130_fd_sc_hd__nor2_1 _21686_ (.A(_04913_),
    .B(_08973_),
    .Y(_01360_));
 sky130_fd_sc_hd__nor2_1 _21687_ (.A(_04923_),
    .B(_08973_),
    .Y(_01361_));
 sky130_fd_sc_hd__nor2_1 _21688_ (.A(_04932_),
    .B(_08973_),
    .Y(_01362_));
 sky130_fd_sc_hd__nor2_1 _21689_ (.A(_04939_),
    .B(_08973_),
    .Y(_01363_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_825 ();
 sky130_fd_sc_hd__nor2_1 _21691_ (.A(_04951_),
    .B(_08973_),
    .Y(_01364_));
 sky130_fd_sc_hd__nor2_1 _21692_ (.A(_04794_),
    .B(_08973_),
    .Y(_01365_));
 sky130_fd_sc_hd__nor2_1 _21693_ (.A(_04960_),
    .B(_08973_),
    .Y(_01366_));
 sky130_fd_sc_hd__nor2_1 _21694_ (.A(_04974_),
    .B(_08973_),
    .Y(_01367_));
 sky130_fd_sc_hd__nor2_1 _21695_ (.A(net1137),
    .B(_08973_),
    .Y(_01368_));
 sky130_fd_sc_hd__nor2_1 _21696_ (.A(_04990_),
    .B(_08973_),
    .Y(_01369_));
 sky130_fd_sc_hd__nor2_1 _21697_ (.A(net1128),
    .B(_08973_),
    .Y(_01370_));
 sky130_fd_sc_hd__nor2_1 _21698_ (.A(_05011_),
    .B(_08973_),
    .Y(_01371_));
 sky130_fd_sc_hd__nor2_1 _21699_ (.A(net1139),
    .B(_08973_),
    .Y(_01372_));
 sky130_fd_sc_hd__nor2_1 _21700_ (.A(_05029_),
    .B(_08973_),
    .Y(_01373_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_824 ();
 sky130_fd_sc_hd__nor2_1 _21702_ (.A(net1135),
    .B(_08973_),
    .Y(_01374_));
 sky130_fd_sc_hd__nor2_1 _21703_ (.A(_05044_),
    .B(_08973_),
    .Y(_01375_));
 sky130_fd_sc_hd__nor2_1 _21704_ (.A(_04801_),
    .B(_08973_),
    .Y(_01376_));
 sky130_fd_sc_hd__nor2_1 _21705_ (.A(_05060_),
    .B(_08973_),
    .Y(_01377_));
 sky130_fd_sc_hd__nor2_1 _21706_ (.A(_08895_),
    .B(_08973_),
    .Y(_01378_));
 sky130_fd_sc_hd__nor2_1 _21707_ (.A(_04808_),
    .B(_08973_),
    .Y(_01379_));
 sky130_fd_sc_hd__nor2_1 _21708_ (.A(_04817_),
    .B(_08973_),
    .Y(_01380_));
 sky130_fd_sc_hd__nor2_1 _21709_ (.A(_04826_),
    .B(_08973_),
    .Y(_01381_));
 sky130_fd_sc_hd__nor2_1 _21710_ (.A(_04834_),
    .B(_08973_),
    .Y(_01382_));
 sky130_fd_sc_hd__nor2_1 _21711_ (.A(_04843_),
    .B(_08973_),
    .Y(_01383_));
 sky130_fd_sc_hd__nor2_1 _21712_ (.A(_04852_),
    .B(_08973_),
    .Y(_01384_));
 sky130_fd_sc_hd__nor2_1 _21713_ (.A(_04860_),
    .B(_08973_),
    .Y(_01385_));
 sky130_fd_sc_hd__nand2_8 _21714_ (.A(_09805_),
    .B(_05474_),
    .Y(_08977_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_823 ();
 sky130_fd_sc_hd__nor2_1 _21716_ (.A(_05118_),
    .B(_08977_),
    .Y(_01386_));
 sky130_fd_sc_hd__nor2_1 _21717_ (.A(_05192_),
    .B(_08977_),
    .Y(_01387_));
 sky130_fd_sc_hd__nor2_1 _21718_ (.A(_05204_),
    .B(_08977_),
    .Y(_01388_));
 sky130_fd_sc_hd__nor2_1 _21719_ (.A(_05214_),
    .B(_08977_),
    .Y(_01389_));
 sky130_fd_sc_hd__nor2_1 _21720_ (.A(_05221_),
    .B(_08977_),
    .Y(_01390_));
 sky130_fd_sc_hd__nor2_1 _21721_ (.A(net1138),
    .B(_08977_),
    .Y(_01391_));
 sky130_fd_sc_hd__nor2_1 _21722_ (.A(_05238_),
    .B(_08977_),
    .Y(_01392_));
 sky130_fd_sc_hd__nor2_1 _21723_ (.A(net1140),
    .B(_08977_),
    .Y(_01393_));
 sky130_fd_sc_hd__nor2_1 _21724_ (.A(_05258_),
    .B(_08977_),
    .Y(_01394_));
 sky130_fd_sc_hd__nor2_1 _21725_ (.A(_05267_),
    .B(_08977_),
    .Y(_01395_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_822 ();
 sky130_fd_sc_hd__nor2_1 _21727_ (.A(_05280_),
    .B(_08977_),
    .Y(_01396_));
 sky130_fd_sc_hd__nor2_1 _21728_ (.A(_05122_),
    .B(_08977_),
    .Y(_01397_));
 sky130_fd_sc_hd__nor2_1 _21729_ (.A(_05291_),
    .B(_08977_),
    .Y(_01398_));
 sky130_fd_sc_hd__nor2_1 _21730_ (.A(_05301_),
    .B(_08977_),
    .Y(_01399_));
 sky130_fd_sc_hd__nor2_1 _21731_ (.A(_05309_),
    .B(_08977_),
    .Y(_01400_));
 sky130_fd_sc_hd__nor2_1 _21732_ (.A(_05320_),
    .B(_08977_),
    .Y(_01401_));
 sky130_fd_sc_hd__nor2_1 _21733_ (.A(net1145),
    .B(_08977_),
    .Y(_01402_));
 sky130_fd_sc_hd__nor2_1 _21734_ (.A(_05339_),
    .B(_08977_),
    .Y(_01403_));
 sky130_fd_sc_hd__nor2_1 _21735_ (.A(net1144),
    .B(_08977_),
    .Y(_01404_));
 sky130_fd_sc_hd__nor2_1 _21736_ (.A(_05358_),
    .B(_08977_),
    .Y(_01405_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_821 ();
 sky130_fd_sc_hd__nor2_1 _21738_ (.A(net1141),
    .B(_08977_),
    .Y(_01406_));
 sky130_fd_sc_hd__nor2_1 _21739_ (.A(_05380_),
    .B(_08977_),
    .Y(_01407_));
 sky130_fd_sc_hd__nor2_1 _21740_ (.A(_05126_),
    .B(_08977_),
    .Y(_01408_));
 sky130_fd_sc_hd__nor2_1 _21741_ (.A(net1114),
    .B(_08977_),
    .Y(_01409_));
 sky130_fd_sc_hd__nor2_1 _21742_ (.A(_05430_),
    .B(_08977_),
    .Y(_01410_));
 sky130_fd_sc_hd__nor2_1 _21743_ (.A(_05132_),
    .B(_08977_),
    .Y(_01411_));
 sky130_fd_sc_hd__nor2_1 _21744_ (.A(_05140_),
    .B(_08977_),
    .Y(_01412_));
 sky130_fd_sc_hd__nor2_1 _21745_ (.A(_05149_),
    .B(_08977_),
    .Y(_01413_));
 sky130_fd_sc_hd__nor2_1 _21746_ (.A(_05157_),
    .B(_08977_),
    .Y(_01414_));
 sky130_fd_sc_hd__nor2_1 _21747_ (.A(_05166_),
    .B(_08977_),
    .Y(_01415_));
 sky130_fd_sc_hd__nor2_1 _21748_ (.A(_05173_),
    .B(_08977_),
    .Y(_01416_));
 sky130_fd_sc_hd__nor2_1 _21749_ (.A(_05183_),
    .B(_08977_),
    .Y(_01417_));
 sky130_fd_sc_hd__nand2_8 _21750_ (.A(_09751_),
    .B(_05516_),
    .Y(_08981_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_820 ();
 sky130_fd_sc_hd__nor2_1 _21752_ (.A(_04790_),
    .B(_08981_),
    .Y(_01418_));
 sky130_fd_sc_hd__nor2_1 _21753_ (.A(_04871_),
    .B(_08981_),
    .Y(_01419_));
 sky130_fd_sc_hd__nor2_1 _21754_ (.A(_04883_),
    .B(_08981_),
    .Y(_01420_));
 sky130_fd_sc_hd__nor2_1 _21755_ (.A(_04892_),
    .B(_08981_),
    .Y(_01421_));
 sky130_fd_sc_hd__nor2_1 _21756_ (.A(_04899_),
    .B(_08981_),
    .Y(_01422_));
 sky130_fd_sc_hd__nor2_1 _21757_ (.A(_04906_),
    .B(_08981_),
    .Y(_01423_));
 sky130_fd_sc_hd__nor2_1 _21758_ (.A(_04913_),
    .B(_08981_),
    .Y(_01424_));
 sky130_fd_sc_hd__nor2_1 _21759_ (.A(_04923_),
    .B(_08981_),
    .Y(_01425_));
 sky130_fd_sc_hd__nor2_1 _21760_ (.A(_04932_),
    .B(_08981_),
    .Y(_01426_));
 sky130_fd_sc_hd__nor2_1 _21761_ (.A(_04939_),
    .B(_08981_),
    .Y(_01427_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_819 ();
 sky130_fd_sc_hd__nor2_1 _21763_ (.A(_04951_),
    .B(_08981_),
    .Y(_01428_));
 sky130_fd_sc_hd__nor2_1 _21764_ (.A(_04794_),
    .B(_08981_),
    .Y(_01429_));
 sky130_fd_sc_hd__nor2_1 _21765_ (.A(_04960_),
    .B(_08981_),
    .Y(_01430_));
 sky130_fd_sc_hd__nor2_1 _21766_ (.A(_04974_),
    .B(_08981_),
    .Y(_01431_));
 sky130_fd_sc_hd__nor2_1 _21767_ (.A(net1137),
    .B(_08981_),
    .Y(_01432_));
 sky130_fd_sc_hd__nor2_1 _21768_ (.A(_04990_),
    .B(_08981_),
    .Y(_01433_));
 sky130_fd_sc_hd__nor2_1 _21769_ (.A(net1128),
    .B(_08981_),
    .Y(_01434_));
 sky130_fd_sc_hd__nor2_1 _21770_ (.A(_05011_),
    .B(_08981_),
    .Y(_01435_));
 sky130_fd_sc_hd__nor2_1 _21771_ (.A(net1139),
    .B(_08981_),
    .Y(_01436_));
 sky130_fd_sc_hd__nor2_1 _21772_ (.A(_05029_),
    .B(_08981_),
    .Y(_01437_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_818 ();
 sky130_fd_sc_hd__nor2_1 _21774_ (.A(_05035_),
    .B(_08981_),
    .Y(_01438_));
 sky130_fd_sc_hd__nor2_1 _21775_ (.A(_05044_),
    .B(_08981_),
    .Y(_01439_));
 sky130_fd_sc_hd__nor2_1 _21776_ (.A(_04801_),
    .B(_08981_),
    .Y(_01440_));
 sky130_fd_sc_hd__nor2_1 _21777_ (.A(_05060_),
    .B(_08981_),
    .Y(_01441_));
 sky130_fd_sc_hd__nor2_1 _21778_ (.A(_08895_),
    .B(_08981_),
    .Y(_01442_));
 sky130_fd_sc_hd__nor2_1 _21779_ (.A(_04808_),
    .B(_08981_),
    .Y(_01443_));
 sky130_fd_sc_hd__nor2_1 _21780_ (.A(_04817_),
    .B(_08981_),
    .Y(_01444_));
 sky130_fd_sc_hd__nor2_1 _21781_ (.A(_04826_),
    .B(_08981_),
    .Y(_01445_));
 sky130_fd_sc_hd__nor2_1 _21782_ (.A(_04834_),
    .B(_08981_),
    .Y(_01446_));
 sky130_fd_sc_hd__nor2_1 _21783_ (.A(_04843_),
    .B(_08981_),
    .Y(_01447_));
 sky130_fd_sc_hd__nor2_1 _21784_ (.A(_04852_),
    .B(_08981_),
    .Y(_01448_));
 sky130_fd_sc_hd__nor2_1 _21785_ (.A(_04860_),
    .B(_08981_),
    .Y(_01449_));
 sky130_fd_sc_hd__nand2_8 _21786_ (.A(_09805_),
    .B(_05557_),
    .Y(_08985_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_817 ();
 sky130_fd_sc_hd__nor2_1 _21788_ (.A(_05118_),
    .B(_08985_),
    .Y(_01450_));
 sky130_fd_sc_hd__nor2_1 _21789_ (.A(_05192_),
    .B(_08985_),
    .Y(_01451_));
 sky130_fd_sc_hd__nor2_1 _21790_ (.A(_05204_),
    .B(_08985_),
    .Y(_01452_));
 sky130_fd_sc_hd__nor2_1 _21791_ (.A(_05214_),
    .B(_08985_),
    .Y(_01453_));
 sky130_fd_sc_hd__nor2_1 _21792_ (.A(_05221_),
    .B(_08985_),
    .Y(_01454_));
 sky130_fd_sc_hd__nor2_1 _21793_ (.A(net1138),
    .B(_08985_),
    .Y(_01455_));
 sky130_fd_sc_hd__nor2_1 _21794_ (.A(_05238_),
    .B(_08985_),
    .Y(_01456_));
 sky130_fd_sc_hd__nor2_1 _21795_ (.A(net1140),
    .B(_08985_),
    .Y(_01457_));
 sky130_fd_sc_hd__nor2_1 _21796_ (.A(_05258_),
    .B(_08985_),
    .Y(_01458_));
 sky130_fd_sc_hd__nor2_1 _21797_ (.A(net1136),
    .B(_08985_),
    .Y(_01459_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_816 ();
 sky130_fd_sc_hd__nor2_1 _21799_ (.A(_05280_),
    .B(_08985_),
    .Y(_01460_));
 sky130_fd_sc_hd__nor2_1 _21800_ (.A(_05122_),
    .B(_08985_),
    .Y(_01461_));
 sky130_fd_sc_hd__nor2_1 _21801_ (.A(_05291_),
    .B(_08985_),
    .Y(_01462_));
 sky130_fd_sc_hd__nor2_1 _21802_ (.A(_05301_),
    .B(_08985_),
    .Y(_01463_));
 sky130_fd_sc_hd__nor2_1 _21803_ (.A(_05309_),
    .B(_08985_),
    .Y(_01464_));
 sky130_fd_sc_hd__nor2_1 _21804_ (.A(_05320_),
    .B(_08985_),
    .Y(_01465_));
 sky130_fd_sc_hd__nor2_1 _21805_ (.A(net1145),
    .B(_08985_),
    .Y(_01466_));
 sky130_fd_sc_hd__nor2_1 _21806_ (.A(_05339_),
    .B(_08985_),
    .Y(_01467_));
 sky130_fd_sc_hd__nor2_1 _21807_ (.A(net1144),
    .B(_08985_),
    .Y(_01468_));
 sky130_fd_sc_hd__nor2_1 _21808_ (.A(_05358_),
    .B(_08985_),
    .Y(_01469_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_815 ();
 sky130_fd_sc_hd__nor2_1 _21810_ (.A(net1134),
    .B(_08985_),
    .Y(_01470_));
 sky130_fd_sc_hd__nor2_1 _21811_ (.A(_05380_),
    .B(_08985_),
    .Y(_01471_));
 sky130_fd_sc_hd__nor2_1 _21812_ (.A(_05126_),
    .B(_08985_),
    .Y(_01472_));
 sky130_fd_sc_hd__nor2_1 _21813_ (.A(net1143),
    .B(_08985_),
    .Y(_01473_));
 sky130_fd_sc_hd__nor2_1 _21814_ (.A(_05430_),
    .B(_08985_),
    .Y(_01474_));
 sky130_fd_sc_hd__nor2_1 _21815_ (.A(_05132_),
    .B(_08985_),
    .Y(_01475_));
 sky130_fd_sc_hd__nor2_1 _21816_ (.A(_05140_),
    .B(_08985_),
    .Y(_01476_));
 sky130_fd_sc_hd__nor2_1 _21817_ (.A(_05149_),
    .B(_08985_),
    .Y(_01477_));
 sky130_fd_sc_hd__nor2_1 _21818_ (.A(_05157_),
    .B(_08985_),
    .Y(_01478_));
 sky130_fd_sc_hd__nor2_1 _21819_ (.A(_05166_),
    .B(_08985_),
    .Y(_01479_));
 sky130_fd_sc_hd__nor2_1 _21820_ (.A(_05173_),
    .B(_08985_),
    .Y(_01480_));
 sky130_fd_sc_hd__nor2_1 _21821_ (.A(_05183_),
    .B(_08985_),
    .Y(_01481_));
 sky130_fd_sc_hd__nand2_8 _21822_ (.A(_09751_),
    .B(_05598_),
    .Y(_08989_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_814 ();
 sky130_fd_sc_hd__nor2_1 _21824_ (.A(_04790_),
    .B(_08989_),
    .Y(_01482_));
 sky130_fd_sc_hd__nor2_1 _21825_ (.A(_04871_),
    .B(_08989_),
    .Y(_01483_));
 sky130_fd_sc_hd__nor2_1 _21826_ (.A(_04883_),
    .B(_08989_),
    .Y(_01484_));
 sky130_fd_sc_hd__nor2_1 _21827_ (.A(_04892_),
    .B(_08989_),
    .Y(_01485_));
 sky130_fd_sc_hd__nor2_1 _21828_ (.A(_04899_),
    .B(_08989_),
    .Y(_01486_));
 sky130_fd_sc_hd__nor2_1 _21829_ (.A(_04906_),
    .B(_08989_),
    .Y(_01487_));
 sky130_fd_sc_hd__nor2_1 _21830_ (.A(_04913_),
    .B(_08989_),
    .Y(_01488_));
 sky130_fd_sc_hd__nor2_1 _21831_ (.A(_04923_),
    .B(_08989_),
    .Y(_01489_));
 sky130_fd_sc_hd__nor2_1 _21832_ (.A(_04932_),
    .B(_08989_),
    .Y(_01490_));
 sky130_fd_sc_hd__nor2_1 _21833_ (.A(_04939_),
    .B(_08989_),
    .Y(_01491_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_813 ();
 sky130_fd_sc_hd__nor2_1 _21835_ (.A(_04951_),
    .B(_08989_),
    .Y(_01492_));
 sky130_fd_sc_hd__nor2_1 _21836_ (.A(_04794_),
    .B(_08989_),
    .Y(_01493_));
 sky130_fd_sc_hd__nor2_1 _21837_ (.A(_04960_),
    .B(_08989_),
    .Y(_01494_));
 sky130_fd_sc_hd__nor2_1 _21838_ (.A(_04974_),
    .B(_08989_),
    .Y(_01495_));
 sky130_fd_sc_hd__nor2_1 _21839_ (.A(net1137),
    .B(_08989_),
    .Y(_01496_));
 sky130_fd_sc_hd__nor2_1 _21840_ (.A(_04990_),
    .B(_08989_),
    .Y(_01497_));
 sky130_fd_sc_hd__nor2_1 _21841_ (.A(net1129),
    .B(_08989_),
    .Y(_01498_));
 sky130_fd_sc_hd__nor2_1 _21842_ (.A(_05011_),
    .B(_08989_),
    .Y(_01499_));
 sky130_fd_sc_hd__nor2_1 _21843_ (.A(_05020_),
    .B(_08989_),
    .Y(_01500_));
 sky130_fd_sc_hd__nor2_1 _21844_ (.A(_05029_),
    .B(_08989_),
    .Y(_01501_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_812 ();
 sky130_fd_sc_hd__nor2_1 _21846_ (.A(net1135),
    .B(_08989_),
    .Y(_01502_));
 sky130_fd_sc_hd__nor2_1 _21847_ (.A(_05044_),
    .B(_08989_),
    .Y(_01503_));
 sky130_fd_sc_hd__nor2_1 _21848_ (.A(_04801_),
    .B(_08989_),
    .Y(_01504_));
 sky130_fd_sc_hd__nor2_1 _21849_ (.A(_05060_),
    .B(_08989_),
    .Y(_01505_));
 sky130_fd_sc_hd__nor2_1 _21850_ (.A(_08895_),
    .B(_08989_),
    .Y(_01506_));
 sky130_fd_sc_hd__nor2_1 _21851_ (.A(_04808_),
    .B(_08989_),
    .Y(_01507_));
 sky130_fd_sc_hd__nor2_1 _21852_ (.A(_04817_),
    .B(_08989_),
    .Y(_01508_));
 sky130_fd_sc_hd__nor2_1 _21853_ (.A(_04826_),
    .B(_08989_),
    .Y(_01509_));
 sky130_fd_sc_hd__nor2_1 _21854_ (.A(_04834_),
    .B(_08989_),
    .Y(_01510_));
 sky130_fd_sc_hd__nor2_1 _21855_ (.A(_04843_),
    .B(_08989_),
    .Y(_01511_));
 sky130_fd_sc_hd__nor2_1 _21856_ (.A(_04852_),
    .B(_08989_),
    .Y(_01512_));
 sky130_fd_sc_hd__nor2_1 _21857_ (.A(_04860_),
    .B(_08989_),
    .Y(_01513_));
 sky130_fd_sc_hd__nand2_8 _21858_ (.A(_09805_),
    .B(_05951_),
    .Y(_08993_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_811 ();
 sky130_fd_sc_hd__nor2_1 _21860_ (.A(_05118_),
    .B(_08993_),
    .Y(_01514_));
 sky130_fd_sc_hd__nor2_1 _21861_ (.A(_05192_),
    .B(_08993_),
    .Y(_01515_));
 sky130_fd_sc_hd__nor2_1 _21862_ (.A(_05204_),
    .B(_08993_),
    .Y(_01516_));
 sky130_fd_sc_hd__nor2_1 _21863_ (.A(_05214_),
    .B(_08993_),
    .Y(_01517_));
 sky130_fd_sc_hd__nor2_1 _21864_ (.A(_05221_),
    .B(_08993_),
    .Y(_01518_));
 sky130_fd_sc_hd__nor2_1 _21865_ (.A(_05228_),
    .B(_08993_),
    .Y(_01519_));
 sky130_fd_sc_hd__nor2_1 _21866_ (.A(_05238_),
    .B(_08993_),
    .Y(_01520_));
 sky130_fd_sc_hd__nor2_1 _21867_ (.A(_05247_),
    .B(_08993_),
    .Y(_01521_));
 sky130_fd_sc_hd__nor2_1 _21868_ (.A(_05258_),
    .B(_08993_),
    .Y(_01522_));
 sky130_fd_sc_hd__nor2_1 _21869_ (.A(net1136),
    .B(_08993_),
    .Y(_01523_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_810 ();
 sky130_fd_sc_hd__nor2_1 _21871_ (.A(_05280_),
    .B(_08993_),
    .Y(_01524_));
 sky130_fd_sc_hd__nor2_1 _21872_ (.A(_05122_),
    .B(_08993_),
    .Y(_01525_));
 sky130_fd_sc_hd__nor2_1 _21873_ (.A(_05291_),
    .B(_08993_),
    .Y(_01526_));
 sky130_fd_sc_hd__nor2_1 _21874_ (.A(_05301_),
    .B(_08993_),
    .Y(_01527_));
 sky130_fd_sc_hd__nor2_1 _21875_ (.A(_05309_),
    .B(_08993_),
    .Y(_01528_));
 sky130_fd_sc_hd__nor2_1 _21876_ (.A(_05320_),
    .B(_08993_),
    .Y(_01529_));
 sky130_fd_sc_hd__nor2_1 _21877_ (.A(net1145),
    .B(_08993_),
    .Y(_01530_));
 sky130_fd_sc_hd__nor2_1 _21878_ (.A(_05339_),
    .B(_08993_),
    .Y(_01531_));
 sky130_fd_sc_hd__nor2_1 _21879_ (.A(_05347_),
    .B(_08993_),
    .Y(_01532_));
 sky130_fd_sc_hd__nor2_1 _21880_ (.A(_05358_),
    .B(_08993_),
    .Y(_01533_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_809 ();
 sky130_fd_sc_hd__nor2_1 _21882_ (.A(net1134),
    .B(_08993_),
    .Y(_01534_));
 sky130_fd_sc_hd__nor2_1 _21883_ (.A(_05380_),
    .B(_08993_),
    .Y(_01535_));
 sky130_fd_sc_hd__nor2_1 _21884_ (.A(_05126_),
    .B(_08993_),
    .Y(_01536_));
 sky130_fd_sc_hd__nor2_1 _21885_ (.A(net1114),
    .B(_08993_),
    .Y(_01537_));
 sky130_fd_sc_hd__nor2_1 _21886_ (.A(_05430_),
    .B(_08993_),
    .Y(_01538_));
 sky130_fd_sc_hd__nor2_1 _21887_ (.A(_05132_),
    .B(_08993_),
    .Y(_01539_));
 sky130_fd_sc_hd__nor2_1 _21888_ (.A(_05140_),
    .B(_08993_),
    .Y(_01540_));
 sky130_fd_sc_hd__nor2_1 _21889_ (.A(_05149_),
    .B(_08993_),
    .Y(_01541_));
 sky130_fd_sc_hd__nor2_1 _21890_ (.A(_05157_),
    .B(_08993_),
    .Y(_01542_));
 sky130_fd_sc_hd__nor2_1 _21891_ (.A(_05166_),
    .B(_08993_),
    .Y(_01543_));
 sky130_fd_sc_hd__nor2_1 _21892_ (.A(_05173_),
    .B(_08993_),
    .Y(_01544_));
 sky130_fd_sc_hd__nor2_1 _21893_ (.A(_05183_),
    .B(_08993_),
    .Y(_01545_));
 sky130_fd_sc_hd__nand2_8 _21894_ (.A(_09759_),
    .B(_04784_),
    .Y(_08997_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_808 ();
 sky130_fd_sc_hd__nor2_1 _21896_ (.A(_04790_),
    .B(_08997_),
    .Y(_01546_));
 sky130_fd_sc_hd__nor2_1 _21897_ (.A(_04871_),
    .B(_08997_),
    .Y(_01547_));
 sky130_fd_sc_hd__nor2_1 _21898_ (.A(_04883_),
    .B(_08997_),
    .Y(_01548_));
 sky130_fd_sc_hd__nor2_1 _21899_ (.A(_04892_),
    .B(_08997_),
    .Y(_01549_));
 sky130_fd_sc_hd__nor2_1 _21900_ (.A(_04899_),
    .B(_08997_),
    .Y(_01550_));
 sky130_fd_sc_hd__nor2_1 _21901_ (.A(_04906_),
    .B(_08997_),
    .Y(_01551_));
 sky130_fd_sc_hd__nor2_1 _21902_ (.A(_04913_),
    .B(_08997_),
    .Y(_01552_));
 sky130_fd_sc_hd__nor2_1 _21903_ (.A(_04923_),
    .B(_08997_),
    .Y(_01553_));
 sky130_fd_sc_hd__nor2_1 _21904_ (.A(_04932_),
    .B(_08997_),
    .Y(_01554_));
 sky130_fd_sc_hd__nor2_1 _21905_ (.A(net1142),
    .B(_08997_),
    .Y(_01555_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_807 ();
 sky130_fd_sc_hd__nor2_1 _21907_ (.A(_04951_),
    .B(_08997_),
    .Y(_01556_));
 sky130_fd_sc_hd__nor2_1 _21908_ (.A(_04794_),
    .B(_08997_),
    .Y(_01557_));
 sky130_fd_sc_hd__nor2_1 _21909_ (.A(_04960_),
    .B(_08997_),
    .Y(_01558_));
 sky130_fd_sc_hd__nor2_1 _21910_ (.A(_04974_),
    .B(_08997_),
    .Y(_01559_));
 sky130_fd_sc_hd__nor2_1 _21911_ (.A(net1137),
    .B(_08997_),
    .Y(_01560_));
 sky130_fd_sc_hd__nor2_1 _21912_ (.A(_04990_),
    .B(_08997_),
    .Y(_01561_));
 sky130_fd_sc_hd__nor2_1 _21913_ (.A(_05000_),
    .B(_08997_),
    .Y(_01562_));
 sky130_fd_sc_hd__nor2_1 _21914_ (.A(_05011_),
    .B(_08997_),
    .Y(_01563_));
 sky130_fd_sc_hd__nor2_1 _21915_ (.A(_05020_),
    .B(_08997_),
    .Y(_01564_));
 sky130_fd_sc_hd__nor2_1 _21916_ (.A(_05029_),
    .B(_08997_),
    .Y(_01565_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_806 ();
 sky130_fd_sc_hd__nor2_1 _21918_ (.A(_05035_),
    .B(_08997_),
    .Y(_01566_));
 sky130_fd_sc_hd__nor2_1 _21919_ (.A(_05044_),
    .B(_08997_),
    .Y(_01567_));
 sky130_fd_sc_hd__nor2_1 _21920_ (.A(_04801_),
    .B(_08997_),
    .Y(_01568_));
 sky130_fd_sc_hd__nor2_1 _21921_ (.A(_05060_),
    .B(_08997_),
    .Y(_01569_));
 sky130_fd_sc_hd__nor2_1 _21922_ (.A(_08895_),
    .B(_08997_),
    .Y(_01570_));
 sky130_fd_sc_hd__nor2_1 _21923_ (.A(_04808_),
    .B(_08997_),
    .Y(_01571_));
 sky130_fd_sc_hd__nor2_1 _21924_ (.A(_04817_),
    .B(_08997_),
    .Y(_01572_));
 sky130_fd_sc_hd__nor2_1 _21925_ (.A(_04826_),
    .B(_08997_),
    .Y(_01573_));
 sky130_fd_sc_hd__nor2_1 _21926_ (.A(_04834_),
    .B(_08997_),
    .Y(_01574_));
 sky130_fd_sc_hd__nor2_1 _21927_ (.A(_04843_),
    .B(_08997_),
    .Y(_01575_));
 sky130_fd_sc_hd__nor2_1 _21928_ (.A(_04852_),
    .B(_08997_),
    .Y(_01576_));
 sky130_fd_sc_hd__nor2_1 _21929_ (.A(_04860_),
    .B(_08997_),
    .Y(_01577_));
 sky130_fd_sc_hd__nand2_8 _21930_ (.A(_09811_),
    .B(_05115_),
    .Y(_09001_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_805 ();
 sky130_fd_sc_hd__nor2_1 _21932_ (.A(_05118_),
    .B(_09001_),
    .Y(_01578_));
 sky130_fd_sc_hd__nor2_1 _21933_ (.A(_05192_),
    .B(_09001_),
    .Y(_01579_));
 sky130_fd_sc_hd__nor2_1 _21934_ (.A(_05204_),
    .B(_09001_),
    .Y(_01580_));
 sky130_fd_sc_hd__nor2_1 _21935_ (.A(_05214_),
    .B(_09001_),
    .Y(_01581_));
 sky130_fd_sc_hd__nor2_1 _21936_ (.A(_05221_),
    .B(_09001_),
    .Y(_01582_));
 sky130_fd_sc_hd__nor2_1 _21937_ (.A(net1138),
    .B(_09001_),
    .Y(_01583_));
 sky130_fd_sc_hd__nor2_1 _21938_ (.A(_05238_),
    .B(_09001_),
    .Y(_01584_));
 sky130_fd_sc_hd__nor2_1 _21939_ (.A(net1140),
    .B(_09001_),
    .Y(_01585_));
 sky130_fd_sc_hd__nor2_1 _21940_ (.A(_05258_),
    .B(_09001_),
    .Y(_01586_));
 sky130_fd_sc_hd__nor2_1 _21941_ (.A(net1136),
    .B(_09001_),
    .Y(_01587_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_804 ();
 sky130_fd_sc_hd__nor2_1 _21943_ (.A(_05280_),
    .B(_09001_),
    .Y(_01588_));
 sky130_fd_sc_hd__nor2_1 _21944_ (.A(_05122_),
    .B(_09001_),
    .Y(_01589_));
 sky130_fd_sc_hd__nor2_1 _21945_ (.A(_05291_),
    .B(_09001_),
    .Y(_01590_));
 sky130_fd_sc_hd__nor2_1 _21946_ (.A(_05301_),
    .B(_09001_),
    .Y(_01591_));
 sky130_fd_sc_hd__nor2_1 _21947_ (.A(_05309_),
    .B(_09001_),
    .Y(_01592_));
 sky130_fd_sc_hd__nor2_1 _21948_ (.A(_05320_),
    .B(_09001_),
    .Y(_01593_));
 sky130_fd_sc_hd__nor2_1 _21949_ (.A(net1112),
    .B(_09001_),
    .Y(_01594_));
 sky130_fd_sc_hd__nor2_1 _21950_ (.A(_05339_),
    .B(_09001_),
    .Y(_01595_));
 sky130_fd_sc_hd__nor2_1 _21951_ (.A(net1144),
    .B(_09001_),
    .Y(_01596_));
 sky130_fd_sc_hd__nor2_1 _21952_ (.A(_05358_),
    .B(_09001_),
    .Y(_01597_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_803 ();
 sky130_fd_sc_hd__nor2_1 _21954_ (.A(net1141),
    .B(_09001_),
    .Y(_01598_));
 sky130_fd_sc_hd__nor2_1 _21955_ (.A(_05380_),
    .B(_09001_),
    .Y(_01599_));
 sky130_fd_sc_hd__nor2_1 _21956_ (.A(_05126_),
    .B(_09001_),
    .Y(_01600_));
 sky130_fd_sc_hd__nor2_1 _21957_ (.A(net1114),
    .B(_09001_),
    .Y(_01601_));
 sky130_fd_sc_hd__nor2_1 _21958_ (.A(_05430_),
    .B(_09001_),
    .Y(_01602_));
 sky130_fd_sc_hd__nor2_1 _21959_ (.A(_05132_),
    .B(_09001_),
    .Y(_01603_));
 sky130_fd_sc_hd__nor2_1 _21960_ (.A(_05140_),
    .B(_09001_),
    .Y(_01604_));
 sky130_fd_sc_hd__nor2_1 _21961_ (.A(_05149_),
    .B(_09001_),
    .Y(_01605_));
 sky130_fd_sc_hd__nor2_1 _21962_ (.A(_05157_),
    .B(_09001_),
    .Y(_01606_));
 sky130_fd_sc_hd__nor2_1 _21963_ (.A(_05166_),
    .B(_09001_),
    .Y(_01607_));
 sky130_fd_sc_hd__nor2_1 _21964_ (.A(_05173_),
    .B(_09001_),
    .Y(_01608_));
 sky130_fd_sc_hd__nor2_1 _21965_ (.A(_05183_),
    .B(_09001_),
    .Y(_01609_));
 sky130_fd_sc_hd__nand2_8 _21966_ (.A(_09759_),
    .B(_05433_),
    .Y(_09005_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_802 ();
 sky130_fd_sc_hd__nor2_1 _21968_ (.A(_04790_),
    .B(_09005_),
    .Y(_01610_));
 sky130_fd_sc_hd__nor2_1 _21969_ (.A(_04871_),
    .B(_09005_),
    .Y(_01611_));
 sky130_fd_sc_hd__nor2_1 _21970_ (.A(_04883_),
    .B(_09005_),
    .Y(_01612_));
 sky130_fd_sc_hd__nor2_1 _21971_ (.A(_04892_),
    .B(_09005_),
    .Y(_01613_));
 sky130_fd_sc_hd__nor2_1 _21972_ (.A(_04899_),
    .B(_09005_),
    .Y(_01614_));
 sky130_fd_sc_hd__nor2_1 _21973_ (.A(_04906_),
    .B(_09005_),
    .Y(_01615_));
 sky130_fd_sc_hd__nor2_1 _21974_ (.A(_04913_),
    .B(_09005_),
    .Y(_01616_));
 sky130_fd_sc_hd__nor2_1 _21975_ (.A(_04923_),
    .B(_09005_),
    .Y(_01617_));
 sky130_fd_sc_hd__nor2_1 _21976_ (.A(_04932_),
    .B(_09005_),
    .Y(_01618_));
 sky130_fd_sc_hd__nor2_1 _21977_ (.A(net1142),
    .B(_09005_),
    .Y(_01619_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_801 ();
 sky130_fd_sc_hd__nor2_1 _21979_ (.A(_04951_),
    .B(_09005_),
    .Y(_01620_));
 sky130_fd_sc_hd__nor2_1 _21980_ (.A(_04794_),
    .B(_09005_),
    .Y(_01621_));
 sky130_fd_sc_hd__nor2_1 _21981_ (.A(_04960_),
    .B(_09005_),
    .Y(_01622_));
 sky130_fd_sc_hd__nor2_1 _21982_ (.A(_04974_),
    .B(_09005_),
    .Y(_01623_));
 sky130_fd_sc_hd__nor2_1 _21983_ (.A(_04984_),
    .B(_09005_),
    .Y(_01624_));
 sky130_fd_sc_hd__nor2_1 _21984_ (.A(_04990_),
    .B(_09005_),
    .Y(_01625_));
 sky130_fd_sc_hd__nor2_1 _21985_ (.A(net1128),
    .B(_09005_),
    .Y(_01626_));
 sky130_fd_sc_hd__nor2_1 _21986_ (.A(_05011_),
    .B(_09005_),
    .Y(_01627_));
 sky130_fd_sc_hd__nor2_1 _21987_ (.A(net1139),
    .B(_09005_),
    .Y(_01628_));
 sky130_fd_sc_hd__nor2_1 _21988_ (.A(_05029_),
    .B(_09005_),
    .Y(_01629_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_800 ();
 sky130_fd_sc_hd__nor2_1 _21990_ (.A(net1135),
    .B(_09005_),
    .Y(_01630_));
 sky130_fd_sc_hd__nor2_1 _21991_ (.A(_05044_),
    .B(_09005_),
    .Y(_01631_));
 sky130_fd_sc_hd__nor2_1 _21992_ (.A(_04801_),
    .B(_09005_),
    .Y(_01632_));
 sky130_fd_sc_hd__nor2_1 _21993_ (.A(_05060_),
    .B(_09005_),
    .Y(_01633_));
 sky130_fd_sc_hd__nor2_1 _21994_ (.A(_08895_),
    .B(_09005_),
    .Y(_01634_));
 sky130_fd_sc_hd__nor2_1 _21995_ (.A(_04808_),
    .B(_09005_),
    .Y(_01635_));
 sky130_fd_sc_hd__nor2_1 _21996_ (.A(_04817_),
    .B(_09005_),
    .Y(_01636_));
 sky130_fd_sc_hd__nor2_1 _21997_ (.A(_04826_),
    .B(_09005_),
    .Y(_01637_));
 sky130_fd_sc_hd__nor2_1 _21998_ (.A(_04834_),
    .B(_09005_),
    .Y(_01638_));
 sky130_fd_sc_hd__nor2_1 _21999_ (.A(_04843_),
    .B(_09005_),
    .Y(_01639_));
 sky130_fd_sc_hd__nor2_1 _22000_ (.A(_04852_),
    .B(_09005_),
    .Y(_01640_));
 sky130_fd_sc_hd__nor2_1 _22001_ (.A(_04860_),
    .B(_09005_),
    .Y(_01641_));
 sky130_fd_sc_hd__nand2_8 _22002_ (.A(_09811_),
    .B(_05474_),
    .Y(_09009_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_799 ();
 sky130_fd_sc_hd__nor2_1 _22004_ (.A(_05118_),
    .B(_09009_),
    .Y(_01642_));
 sky130_fd_sc_hd__nor2_1 _22005_ (.A(_05192_),
    .B(_09009_),
    .Y(_01643_));
 sky130_fd_sc_hd__nor2_1 _22006_ (.A(_05204_),
    .B(_09009_),
    .Y(_01644_));
 sky130_fd_sc_hd__nor2_1 _22007_ (.A(_05214_),
    .B(_09009_),
    .Y(_01645_));
 sky130_fd_sc_hd__nor2_1 _22008_ (.A(_05221_),
    .B(_09009_),
    .Y(_01646_));
 sky130_fd_sc_hd__nor2_1 _22009_ (.A(_05228_),
    .B(_09009_),
    .Y(_01647_));
 sky130_fd_sc_hd__nor2_1 _22010_ (.A(_05238_),
    .B(_09009_),
    .Y(_01648_));
 sky130_fd_sc_hd__nor2_1 _22011_ (.A(_05247_),
    .B(_09009_),
    .Y(_01649_));
 sky130_fd_sc_hd__nor2_1 _22012_ (.A(_05258_),
    .B(_09009_),
    .Y(_01650_));
 sky130_fd_sc_hd__nor2_1 _22013_ (.A(net1136),
    .B(_09009_),
    .Y(_01651_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_798 ();
 sky130_fd_sc_hd__nor2_1 _22015_ (.A(_05280_),
    .B(_09009_),
    .Y(_01652_));
 sky130_fd_sc_hd__nor2_1 _22016_ (.A(_05122_),
    .B(_09009_),
    .Y(_01653_));
 sky130_fd_sc_hd__nor2_1 _22017_ (.A(_05291_),
    .B(_09009_),
    .Y(_01654_));
 sky130_fd_sc_hd__nor2_1 _22018_ (.A(_05301_),
    .B(_09009_),
    .Y(_01655_));
 sky130_fd_sc_hd__nor2_1 _22019_ (.A(_05309_),
    .B(_09009_),
    .Y(_01656_));
 sky130_fd_sc_hd__nor2_1 _22020_ (.A(_05320_),
    .B(_09009_),
    .Y(_01657_));
 sky130_fd_sc_hd__nor2_1 _22021_ (.A(net1112),
    .B(_09009_),
    .Y(_01658_));
 sky130_fd_sc_hd__nor2_1 _22022_ (.A(_05339_),
    .B(_09009_),
    .Y(_01659_));
 sky130_fd_sc_hd__nor2_1 _22023_ (.A(net1144),
    .B(_09009_),
    .Y(_01660_));
 sky130_fd_sc_hd__nor2_1 _22024_ (.A(_05358_),
    .B(_09009_),
    .Y(_01661_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_797 ();
 sky130_fd_sc_hd__nor2_1 _22026_ (.A(net1141),
    .B(_09009_),
    .Y(_01662_));
 sky130_fd_sc_hd__nor2_1 _22027_ (.A(_05380_),
    .B(_09009_),
    .Y(_01663_));
 sky130_fd_sc_hd__nor2_1 _22028_ (.A(_05126_),
    .B(_09009_),
    .Y(_01664_));
 sky130_fd_sc_hd__nor2_1 _22029_ (.A(net1114),
    .B(_09009_),
    .Y(_01665_));
 sky130_fd_sc_hd__nor2_1 _22030_ (.A(_05430_),
    .B(_09009_),
    .Y(_01666_));
 sky130_fd_sc_hd__nor2_1 _22031_ (.A(_05132_),
    .B(_09009_),
    .Y(_01667_));
 sky130_fd_sc_hd__nor2_1 _22032_ (.A(_05140_),
    .B(_09009_),
    .Y(_01668_));
 sky130_fd_sc_hd__nor2_1 _22033_ (.A(_05149_),
    .B(_09009_),
    .Y(_01669_));
 sky130_fd_sc_hd__nor2_1 _22034_ (.A(_05157_),
    .B(_09009_),
    .Y(_01670_));
 sky130_fd_sc_hd__nor2_1 _22035_ (.A(_05166_),
    .B(_09009_),
    .Y(_01671_));
 sky130_fd_sc_hd__nor2_1 _22036_ (.A(_05173_),
    .B(_09009_),
    .Y(_01672_));
 sky130_fd_sc_hd__nor2_1 _22037_ (.A(_05183_),
    .B(_09009_),
    .Y(_01673_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_796 ();
 sky130_fd_sc_hd__nand2_8 _22039_ (.A(_09759_),
    .B(_05516_),
    .Y(_09014_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_795 ();
 sky130_fd_sc_hd__nor2_1 _22041_ (.A(_04790_),
    .B(_09014_),
    .Y(_01674_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_794 ();
 sky130_fd_sc_hd__nor2_1 _22043_ (.A(_04871_),
    .B(_09014_),
    .Y(_01675_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_793 ();
 sky130_fd_sc_hd__nor2_1 _22045_ (.A(_04883_),
    .B(_09014_),
    .Y(_01676_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_792 ();
 sky130_fd_sc_hd__nor2_1 _22047_ (.A(_04892_),
    .B(_09014_),
    .Y(_01677_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_791 ();
 sky130_fd_sc_hd__nor2_1 _22049_ (.A(_04899_),
    .B(_09014_),
    .Y(_01678_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_790 ();
 sky130_fd_sc_hd__nor2_1 _22051_ (.A(_04906_),
    .B(_09014_),
    .Y(_01679_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_789 ();
 sky130_fd_sc_hd__nor2_1 _22053_ (.A(_04913_),
    .B(_09014_),
    .Y(_01680_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_788 ();
 sky130_fd_sc_hd__nor2_1 _22055_ (.A(_04923_),
    .B(_09014_),
    .Y(_01681_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_787 ();
 sky130_fd_sc_hd__nor2_1 _22057_ (.A(_04932_),
    .B(_09014_),
    .Y(_01682_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_786 ();
 sky130_fd_sc_hd__nor2_1 _22059_ (.A(net1142),
    .B(_09014_),
    .Y(_01683_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_784 ();
 sky130_fd_sc_hd__nor2_1 _22062_ (.A(_04951_),
    .B(_09014_),
    .Y(_01684_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_783 ();
 sky130_fd_sc_hd__nor2_1 _22064_ (.A(_04794_),
    .B(_09014_),
    .Y(_01685_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_782 ();
 sky130_fd_sc_hd__nor2_1 _22066_ (.A(_04960_),
    .B(_09014_),
    .Y(_01686_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_781 ();
 sky130_fd_sc_hd__nor2_1 _22068_ (.A(_04974_),
    .B(_09014_),
    .Y(_01687_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_780 ();
 sky130_fd_sc_hd__nor2_1 _22070_ (.A(_04984_),
    .B(_09014_),
    .Y(_01688_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_779 ();
 sky130_fd_sc_hd__nor2_1 _22072_ (.A(_04990_),
    .B(_09014_),
    .Y(_01689_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_778 ();
 sky130_fd_sc_hd__nor2_1 _22074_ (.A(_05000_),
    .B(_09014_),
    .Y(_01690_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_777 ();
 sky130_fd_sc_hd__nor2_1 _22076_ (.A(_05011_),
    .B(_09014_),
    .Y(_01691_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_776 ();
 sky130_fd_sc_hd__nor2_1 _22078_ (.A(net1139),
    .B(_09014_),
    .Y(_01692_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_775 ();
 sky130_fd_sc_hd__nor2_1 _22080_ (.A(_05029_),
    .B(_09014_),
    .Y(_01693_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_773 ();
 sky130_fd_sc_hd__nor2_1 _22083_ (.A(_05035_),
    .B(_09014_),
    .Y(_01694_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_772 ();
 sky130_fd_sc_hd__nor2_1 _22085_ (.A(_05044_),
    .B(_09014_),
    .Y(_01695_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_771 ();
 sky130_fd_sc_hd__nor2_1 _22087_ (.A(_04801_),
    .B(_09014_),
    .Y(_01696_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_770 ();
 sky130_fd_sc_hd__nor2_1 _22089_ (.A(_05060_),
    .B(_09014_),
    .Y(_01697_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_769 ();
 sky130_fd_sc_hd__nor2_1 _22091_ (.A(_08895_),
    .B(_09014_),
    .Y(_01698_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_768 ();
 sky130_fd_sc_hd__nor2_1 _22093_ (.A(_04808_),
    .B(_09014_),
    .Y(_01699_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_767 ();
 sky130_fd_sc_hd__nor2_1 _22095_ (.A(_04817_),
    .B(_09014_),
    .Y(_01700_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_766 ();
 sky130_fd_sc_hd__nor2_1 _22097_ (.A(_04826_),
    .B(_09014_),
    .Y(_01701_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_765 ();
 sky130_fd_sc_hd__nor2_1 _22099_ (.A(_04834_),
    .B(_09014_),
    .Y(_01702_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_764 ();
 sky130_fd_sc_hd__nor2_1 _22101_ (.A(_04843_),
    .B(_09014_),
    .Y(_01703_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_763 ();
 sky130_fd_sc_hd__nor2_1 _22103_ (.A(_04852_),
    .B(_09014_),
    .Y(_01704_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_762 ();
 sky130_fd_sc_hd__nor2_1 _22105_ (.A(_04860_),
    .B(_09014_),
    .Y(_01705_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_761 ();
 sky130_fd_sc_hd__nand2_8 _22107_ (.A(_09811_),
    .B(_05557_),
    .Y(_09050_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_760 ();
 sky130_fd_sc_hd__nor2_1 _22109_ (.A(_05118_),
    .B(_09050_),
    .Y(_01706_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_759 ();
 sky130_fd_sc_hd__nor2_1 _22111_ (.A(_05192_),
    .B(_09050_),
    .Y(_01707_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_758 ();
 sky130_fd_sc_hd__nor2_1 _22113_ (.A(_05204_),
    .B(_09050_),
    .Y(_01708_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_757 ();
 sky130_fd_sc_hd__nor2_1 _22115_ (.A(_05214_),
    .B(_09050_),
    .Y(_01709_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_756 ();
 sky130_fd_sc_hd__nor2_1 _22117_ (.A(_05221_),
    .B(_09050_),
    .Y(_01710_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_755 ();
 sky130_fd_sc_hd__nor2_1 _22119_ (.A(net1138),
    .B(_09050_),
    .Y(_01711_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_754 ();
 sky130_fd_sc_hd__nor2_1 _22121_ (.A(_05238_),
    .B(_09050_),
    .Y(_01712_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_753 ();
 sky130_fd_sc_hd__nor2_1 _22123_ (.A(net1140),
    .B(_09050_),
    .Y(_01713_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_752 ();
 sky130_fd_sc_hd__nor2_1 _22125_ (.A(_05258_),
    .B(_09050_),
    .Y(_01714_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_751 ();
 sky130_fd_sc_hd__nor2_1 _22127_ (.A(_05267_),
    .B(_09050_),
    .Y(_01715_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_749 ();
 sky130_fd_sc_hd__nor2_1 _22130_ (.A(_05280_),
    .B(_09050_),
    .Y(_01716_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_748 ();
 sky130_fd_sc_hd__nor2_1 _22132_ (.A(_05122_),
    .B(_09050_),
    .Y(_01717_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_747 ();
 sky130_fd_sc_hd__nor2_1 _22134_ (.A(_05291_),
    .B(_09050_),
    .Y(_01718_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_746 ();
 sky130_fd_sc_hd__nor2_1 _22136_ (.A(_05301_),
    .B(_09050_),
    .Y(_01719_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_745 ();
 sky130_fd_sc_hd__nor2_1 _22138_ (.A(_05309_),
    .B(_09050_),
    .Y(_01720_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_744 ();
 sky130_fd_sc_hd__nor2_1 _22140_ (.A(_05320_),
    .B(_09050_),
    .Y(_01721_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_743 ();
 sky130_fd_sc_hd__nor2_1 _22142_ (.A(net1112),
    .B(_09050_),
    .Y(_01722_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_742 ();
 sky130_fd_sc_hd__nor2_1 _22144_ (.A(_05339_),
    .B(_09050_),
    .Y(_01723_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_741 ();
 sky130_fd_sc_hd__nor2_1 _22146_ (.A(net1144),
    .B(_09050_),
    .Y(_01724_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_740 ();
 sky130_fd_sc_hd__nor2_1 _22148_ (.A(_05358_),
    .B(_09050_),
    .Y(_01725_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_738 ();
 sky130_fd_sc_hd__nor2_1 _22151_ (.A(net1113),
    .B(_09050_),
    .Y(_01726_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_737 ();
 sky130_fd_sc_hd__nor2_1 _22153_ (.A(_05380_),
    .B(_09050_),
    .Y(_01727_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_736 ();
 sky130_fd_sc_hd__nor2_1 _22155_ (.A(_05126_),
    .B(_09050_),
    .Y(_01728_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_735 ();
 sky130_fd_sc_hd__nor2_1 _22157_ (.A(net1114),
    .B(_09050_),
    .Y(_01729_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_734 ();
 sky130_fd_sc_hd__nor2_1 _22159_ (.A(_05430_),
    .B(_09050_),
    .Y(_01730_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_733 ();
 sky130_fd_sc_hd__nor2_1 _22161_ (.A(_05132_),
    .B(_09050_),
    .Y(_01731_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_732 ();
 sky130_fd_sc_hd__nor2_1 _22163_ (.A(_05140_),
    .B(_09050_),
    .Y(_01732_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_731 ();
 sky130_fd_sc_hd__nor2_1 _22165_ (.A(_05149_),
    .B(_09050_),
    .Y(_01733_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_730 ();
 sky130_fd_sc_hd__nor2_1 _22167_ (.A(_05157_),
    .B(_09050_),
    .Y(_01734_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_729 ();
 sky130_fd_sc_hd__nor2_1 _22169_ (.A(_05166_),
    .B(_09050_),
    .Y(_01735_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_728 ();
 sky130_fd_sc_hd__nor2_1 _22171_ (.A(_05173_),
    .B(_09050_),
    .Y(_01736_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_727 ();
 sky130_fd_sc_hd__nor2_1 _22173_ (.A(_05183_),
    .B(_09050_),
    .Y(_01737_));
 sky130_fd_sc_hd__nand2_8 _22174_ (.A(_09759_),
    .B(_05598_),
    .Y(_09085_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_726 ();
 sky130_fd_sc_hd__nor2_1 _22176_ (.A(_04790_),
    .B(_09085_),
    .Y(_01738_));
 sky130_fd_sc_hd__nor2_1 _22177_ (.A(_04871_),
    .B(_09085_),
    .Y(_01739_));
 sky130_fd_sc_hd__nor2_1 _22178_ (.A(_04883_),
    .B(_09085_),
    .Y(_01740_));
 sky130_fd_sc_hd__nor2_1 _22179_ (.A(_04892_),
    .B(_09085_),
    .Y(_01741_));
 sky130_fd_sc_hd__nor2_1 _22180_ (.A(_04899_),
    .B(_09085_),
    .Y(_01742_));
 sky130_fd_sc_hd__nor2_1 _22181_ (.A(_04906_),
    .B(_09085_),
    .Y(_01743_));
 sky130_fd_sc_hd__nor2_1 _22182_ (.A(_04913_),
    .B(_09085_),
    .Y(_01744_));
 sky130_fd_sc_hd__nor2_1 _22183_ (.A(_04923_),
    .B(_09085_),
    .Y(_01745_));
 sky130_fd_sc_hd__nor2_1 _22184_ (.A(_04932_),
    .B(_09085_),
    .Y(_01746_));
 sky130_fd_sc_hd__nor2_1 _22185_ (.A(_04939_),
    .B(_09085_),
    .Y(_01747_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_725 ();
 sky130_fd_sc_hd__nor2_1 _22187_ (.A(_04951_),
    .B(_09085_),
    .Y(_01748_));
 sky130_fd_sc_hd__nor2_1 _22188_ (.A(_04794_),
    .B(_09085_),
    .Y(_01749_));
 sky130_fd_sc_hd__nor2_1 _22189_ (.A(_04960_),
    .B(_09085_),
    .Y(_01750_));
 sky130_fd_sc_hd__nor2_1 _22190_ (.A(_04974_),
    .B(_09085_),
    .Y(_01751_));
 sky130_fd_sc_hd__nor2_1 _22191_ (.A(_04984_),
    .B(_09085_),
    .Y(_01752_));
 sky130_fd_sc_hd__nor2_1 _22192_ (.A(_04990_),
    .B(_09085_),
    .Y(_01753_));
 sky130_fd_sc_hd__nor2_1 _22193_ (.A(net1128),
    .B(_09085_),
    .Y(_01754_));
 sky130_fd_sc_hd__nor2_1 _22194_ (.A(_05011_),
    .B(_09085_),
    .Y(_01755_));
 sky130_fd_sc_hd__nor2_1 _22195_ (.A(net1139),
    .B(_09085_),
    .Y(_01756_));
 sky130_fd_sc_hd__nor2_1 _22196_ (.A(_05029_),
    .B(_09085_),
    .Y(_01757_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_724 ();
 sky130_fd_sc_hd__nor2_1 _22198_ (.A(net1135),
    .B(_09085_),
    .Y(_01758_));
 sky130_fd_sc_hd__nor2_1 _22199_ (.A(_05044_),
    .B(_09085_),
    .Y(_01759_));
 sky130_fd_sc_hd__nor2_1 _22200_ (.A(_04801_),
    .B(_09085_),
    .Y(_01760_));
 sky130_fd_sc_hd__nor2_1 _22201_ (.A(_05060_),
    .B(_09085_),
    .Y(_01761_));
 sky130_fd_sc_hd__nor2_1 _22202_ (.A(_08895_),
    .B(_09085_),
    .Y(_01762_));
 sky130_fd_sc_hd__nor2_1 _22203_ (.A(_04808_),
    .B(_09085_),
    .Y(_01763_));
 sky130_fd_sc_hd__nor2_1 _22204_ (.A(_04817_),
    .B(_09085_),
    .Y(_01764_));
 sky130_fd_sc_hd__nor2_1 _22205_ (.A(_04826_),
    .B(_09085_),
    .Y(_01765_));
 sky130_fd_sc_hd__nor2_1 _22206_ (.A(_04834_),
    .B(_09085_),
    .Y(_01766_));
 sky130_fd_sc_hd__nor2_1 _22207_ (.A(_04843_),
    .B(_09085_),
    .Y(_01767_));
 sky130_fd_sc_hd__nor2_1 _22208_ (.A(_04852_),
    .B(_09085_),
    .Y(_01768_));
 sky130_fd_sc_hd__nor2_1 _22209_ (.A(_04860_),
    .B(_09085_),
    .Y(_01769_));
 sky130_fd_sc_hd__or4_4 _22210_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(net1039),
    .D(_09816_),
    .X(_09089_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_722 ();
 sky130_fd_sc_hd__nor2_1 _22213_ (.A(_05118_),
    .B(_09089_),
    .Y(_01770_));
 sky130_fd_sc_hd__nor2_1 _22214_ (.A(_05192_),
    .B(_09089_),
    .Y(_01771_));
 sky130_fd_sc_hd__nor2_1 _22215_ (.A(_05204_),
    .B(_09089_),
    .Y(_01772_));
 sky130_fd_sc_hd__nor2_1 _22216_ (.A(_05214_),
    .B(_09089_),
    .Y(_01773_));
 sky130_fd_sc_hd__nor2_1 _22217_ (.A(_05221_),
    .B(_09089_),
    .Y(_01774_));
 sky130_fd_sc_hd__nor2_1 _22218_ (.A(net1138),
    .B(_09089_),
    .Y(_01775_));
 sky130_fd_sc_hd__nor2_1 _22219_ (.A(_05238_),
    .B(_09089_),
    .Y(_01776_));
 sky130_fd_sc_hd__nor2_1 _22220_ (.A(net1140),
    .B(_09089_),
    .Y(_01777_));
 sky130_fd_sc_hd__nor2_1 _22221_ (.A(_05258_),
    .B(_09089_),
    .Y(_01778_));
 sky130_fd_sc_hd__nor2_1 _22222_ (.A(_05267_),
    .B(_09089_),
    .Y(_01779_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_721 ();
 sky130_fd_sc_hd__nor2_1 _22224_ (.A(_05280_),
    .B(_09089_),
    .Y(_01780_));
 sky130_fd_sc_hd__nor2_1 _22225_ (.A(_05122_),
    .B(_09089_),
    .Y(_01781_));
 sky130_fd_sc_hd__nor2_1 _22226_ (.A(_05291_),
    .B(_09089_),
    .Y(_01782_));
 sky130_fd_sc_hd__nor2_1 _22227_ (.A(_05301_),
    .B(_09089_),
    .Y(_01783_));
 sky130_fd_sc_hd__nor2_1 _22228_ (.A(_05309_),
    .B(_09089_),
    .Y(_01784_));
 sky130_fd_sc_hd__nor2_1 _22229_ (.A(_05320_),
    .B(_09089_),
    .Y(_01785_));
 sky130_fd_sc_hd__nor2_1 _22230_ (.A(net1112),
    .B(_09089_),
    .Y(_01786_));
 sky130_fd_sc_hd__nor2_1 _22231_ (.A(_05339_),
    .B(_09089_),
    .Y(_01787_));
 sky130_fd_sc_hd__nor2_1 _22232_ (.A(net1144),
    .B(_09089_),
    .Y(_01788_));
 sky130_fd_sc_hd__nor2_1 _22233_ (.A(_05358_),
    .B(_09089_),
    .Y(_01789_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_720 ();
 sky130_fd_sc_hd__nor2_1 _22235_ (.A(net1141),
    .B(_09089_),
    .Y(_01790_));
 sky130_fd_sc_hd__nor2_1 _22236_ (.A(_05380_),
    .B(_09089_),
    .Y(_01791_));
 sky130_fd_sc_hd__nor2_1 _22237_ (.A(_05126_),
    .B(_09089_),
    .Y(_01792_));
 sky130_fd_sc_hd__nor2_1 _22238_ (.A(net1114),
    .B(_09089_),
    .Y(_01793_));
 sky130_fd_sc_hd__nor2_1 _22239_ (.A(_05430_),
    .B(_09089_),
    .Y(_01794_));
 sky130_fd_sc_hd__nor2_1 _22240_ (.A(_05132_),
    .B(_09089_),
    .Y(_01795_));
 sky130_fd_sc_hd__nor2_1 _22241_ (.A(_05140_),
    .B(_09089_),
    .Y(_01796_));
 sky130_fd_sc_hd__nor2_1 _22242_ (.A(_05149_),
    .B(_09089_),
    .Y(_01797_));
 sky130_fd_sc_hd__nor2_1 _22243_ (.A(_05157_),
    .B(_09089_),
    .Y(_01798_));
 sky130_fd_sc_hd__nor2_1 _22244_ (.A(_05166_),
    .B(_09089_),
    .Y(_01799_));
 sky130_fd_sc_hd__nor2_1 _22245_ (.A(_05173_),
    .B(_09089_),
    .Y(_01800_));
 sky130_fd_sc_hd__nor2_1 _22246_ (.A(_05183_),
    .B(_09089_),
    .Y(_01801_));
 sky130_fd_sc_hd__nand2_8 _22247_ (.A(_09764_),
    .B(_04784_),
    .Y(_09094_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_719 ();
 sky130_fd_sc_hd__nor2_1 _22249_ (.A(_04790_),
    .B(_09094_),
    .Y(_01802_));
 sky130_fd_sc_hd__nor2_1 _22250_ (.A(_04871_),
    .B(_09094_),
    .Y(_01803_));
 sky130_fd_sc_hd__nor2_1 _22251_ (.A(_04883_),
    .B(_09094_),
    .Y(_01804_));
 sky130_fd_sc_hd__nor2_1 _22252_ (.A(_04892_),
    .B(_09094_),
    .Y(_01805_));
 sky130_fd_sc_hd__nor2_1 _22253_ (.A(_04899_),
    .B(_09094_),
    .Y(_01806_));
 sky130_fd_sc_hd__nor2_1 _22254_ (.A(_04906_),
    .B(_09094_),
    .Y(_01807_));
 sky130_fd_sc_hd__nor2_1 _22255_ (.A(_04913_),
    .B(_09094_),
    .Y(_01808_));
 sky130_fd_sc_hd__nor2_1 _22256_ (.A(_04923_),
    .B(_09094_),
    .Y(_01809_));
 sky130_fd_sc_hd__nor2_1 _22257_ (.A(_04932_),
    .B(_09094_),
    .Y(_01810_));
 sky130_fd_sc_hd__nor2_1 _22258_ (.A(net1142),
    .B(_09094_),
    .Y(_01811_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_718 ();
 sky130_fd_sc_hd__nor2_1 _22260_ (.A(_04951_),
    .B(_09094_),
    .Y(_01812_));
 sky130_fd_sc_hd__nor2_1 _22261_ (.A(_04794_),
    .B(_09094_),
    .Y(_01813_));
 sky130_fd_sc_hd__nor2_1 _22262_ (.A(_04960_),
    .B(_09094_),
    .Y(_01814_));
 sky130_fd_sc_hd__nor2_1 _22263_ (.A(_04974_),
    .B(_09094_),
    .Y(_01815_));
 sky130_fd_sc_hd__nor2_1 _22264_ (.A(net1137),
    .B(_09094_),
    .Y(_01816_));
 sky130_fd_sc_hd__nor2_1 _22265_ (.A(_04990_),
    .B(_09094_),
    .Y(_01817_));
 sky130_fd_sc_hd__nor2_1 _22266_ (.A(net1129),
    .B(_09094_),
    .Y(_01818_));
 sky130_fd_sc_hd__nor2_1 _22267_ (.A(_05011_),
    .B(_09094_),
    .Y(_01819_));
 sky130_fd_sc_hd__nor2_1 _22268_ (.A(net1139),
    .B(_09094_),
    .Y(_01820_));
 sky130_fd_sc_hd__nor2_1 _22269_ (.A(_05029_),
    .B(_09094_),
    .Y(_01821_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_717 ();
 sky130_fd_sc_hd__nor2_1 _22271_ (.A(net1135),
    .B(_09094_),
    .Y(_01822_));
 sky130_fd_sc_hd__nor2_1 _22272_ (.A(_05044_),
    .B(_09094_),
    .Y(_01823_));
 sky130_fd_sc_hd__nor2_1 _22273_ (.A(_04801_),
    .B(_09094_),
    .Y(_01824_));
 sky130_fd_sc_hd__nor2_1 _22274_ (.A(_05060_),
    .B(_09094_),
    .Y(_01825_));
 sky130_fd_sc_hd__nor2_1 _22275_ (.A(_08895_),
    .B(_09094_),
    .Y(_01826_));
 sky130_fd_sc_hd__nor2_1 _22276_ (.A(_04808_),
    .B(_09094_),
    .Y(_01827_));
 sky130_fd_sc_hd__nor2_1 _22277_ (.A(_04817_),
    .B(_09094_),
    .Y(_01828_));
 sky130_fd_sc_hd__nor2_1 _22278_ (.A(_04826_),
    .B(_09094_),
    .Y(_01829_));
 sky130_fd_sc_hd__nor2_1 _22279_ (.A(_04834_),
    .B(_09094_),
    .Y(_01830_));
 sky130_fd_sc_hd__nor2_1 _22280_ (.A(_04843_),
    .B(_09094_),
    .Y(_01831_));
 sky130_fd_sc_hd__nor2_1 _22281_ (.A(_04852_),
    .B(_09094_),
    .Y(_01832_));
 sky130_fd_sc_hd__nor2_1 _22282_ (.A(_04860_),
    .B(_09094_),
    .Y(_01833_));
 sky130_fd_sc_hd__nand2_8 _22283_ (.A(_09818_),
    .B(_05115_),
    .Y(_09098_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_716 ();
 sky130_fd_sc_hd__nor2_1 _22285_ (.A(_05118_),
    .B(_09098_),
    .Y(_01834_));
 sky130_fd_sc_hd__nor2_1 _22286_ (.A(_05192_),
    .B(_09098_),
    .Y(_01835_));
 sky130_fd_sc_hd__nor2_1 _22287_ (.A(_05204_),
    .B(_09098_),
    .Y(_01836_));
 sky130_fd_sc_hd__nor2_1 _22288_ (.A(_05214_),
    .B(_09098_),
    .Y(_01837_));
 sky130_fd_sc_hd__nor2_1 _22289_ (.A(_05221_),
    .B(_09098_),
    .Y(_01838_));
 sky130_fd_sc_hd__nor2_1 _22290_ (.A(net1138),
    .B(_09098_),
    .Y(_01839_));
 sky130_fd_sc_hd__nor2_1 _22291_ (.A(_05238_),
    .B(_09098_),
    .Y(_01840_));
 sky130_fd_sc_hd__nor2_1 _22292_ (.A(net1140),
    .B(_09098_),
    .Y(_01841_));
 sky130_fd_sc_hd__nor2_1 _22293_ (.A(_05258_),
    .B(_09098_),
    .Y(_01842_));
 sky130_fd_sc_hd__nor2_1 _22294_ (.A(_05267_),
    .B(_09098_),
    .Y(_01843_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_715 ();
 sky130_fd_sc_hd__nor2_1 _22296_ (.A(_05280_),
    .B(_09098_),
    .Y(_01844_));
 sky130_fd_sc_hd__nor2_1 _22297_ (.A(_05122_),
    .B(_09098_),
    .Y(_01845_));
 sky130_fd_sc_hd__nor2_1 _22298_ (.A(_05291_),
    .B(_09098_),
    .Y(_01846_));
 sky130_fd_sc_hd__nor2_1 _22299_ (.A(_05301_),
    .B(_09098_),
    .Y(_01847_));
 sky130_fd_sc_hd__nor2_1 _22300_ (.A(_05309_),
    .B(_09098_),
    .Y(_01848_));
 sky130_fd_sc_hd__nor2_1 _22301_ (.A(_05320_),
    .B(_09098_),
    .Y(_01849_));
 sky130_fd_sc_hd__nor2_1 _22302_ (.A(net1112),
    .B(_09098_),
    .Y(_01850_));
 sky130_fd_sc_hd__nor2_1 _22303_ (.A(_05339_),
    .B(_09098_),
    .Y(_01851_));
 sky130_fd_sc_hd__nor2_1 _22304_ (.A(net1144),
    .B(_09098_),
    .Y(_01852_));
 sky130_fd_sc_hd__nor2_1 _22305_ (.A(_05358_),
    .B(_09098_),
    .Y(_01853_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_714 ();
 sky130_fd_sc_hd__nor2_1 _22307_ (.A(net1134),
    .B(_09098_),
    .Y(_01854_));
 sky130_fd_sc_hd__nor2_1 _22308_ (.A(_05380_),
    .B(_09098_),
    .Y(_01855_));
 sky130_fd_sc_hd__nor2_1 _22309_ (.A(_05126_),
    .B(_09098_),
    .Y(_01856_));
 sky130_fd_sc_hd__nor2_1 _22310_ (.A(net1114),
    .B(_09098_),
    .Y(_01857_));
 sky130_fd_sc_hd__nor2_1 _22311_ (.A(_05430_),
    .B(_09098_),
    .Y(_01858_));
 sky130_fd_sc_hd__nor2_1 _22312_ (.A(_05132_),
    .B(_09098_),
    .Y(_01859_));
 sky130_fd_sc_hd__nor2_1 _22313_ (.A(_05140_),
    .B(_09098_),
    .Y(_01860_));
 sky130_fd_sc_hd__nor2_1 _22314_ (.A(_05149_),
    .B(_09098_),
    .Y(_01861_));
 sky130_fd_sc_hd__nor2_1 _22315_ (.A(_05157_),
    .B(_09098_),
    .Y(_01862_));
 sky130_fd_sc_hd__nor2_1 _22316_ (.A(_05166_),
    .B(_09098_),
    .Y(_01863_));
 sky130_fd_sc_hd__nor2_1 _22317_ (.A(_05173_),
    .B(_09098_),
    .Y(_01864_));
 sky130_fd_sc_hd__nor2_1 _22318_ (.A(_05183_),
    .B(_09098_),
    .Y(_01865_));
 sky130_fd_sc_hd__nand2_8 _22319_ (.A(_09764_),
    .B(_05433_),
    .Y(_09102_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_713 ();
 sky130_fd_sc_hd__nor2_1 _22321_ (.A(_04790_),
    .B(_09102_),
    .Y(_01866_));
 sky130_fd_sc_hd__nor2_1 _22322_ (.A(_04871_),
    .B(_09102_),
    .Y(_01867_));
 sky130_fd_sc_hd__nor2_1 _22323_ (.A(_04883_),
    .B(_09102_),
    .Y(_01868_));
 sky130_fd_sc_hd__nor2_1 _22324_ (.A(_04892_),
    .B(_09102_),
    .Y(_01869_));
 sky130_fd_sc_hd__nor2_1 _22325_ (.A(_04899_),
    .B(_09102_),
    .Y(_01870_));
 sky130_fd_sc_hd__nor2_1 _22326_ (.A(_04906_),
    .B(_09102_),
    .Y(_01871_));
 sky130_fd_sc_hd__nor2_1 _22327_ (.A(_04913_),
    .B(_09102_),
    .Y(_01872_));
 sky130_fd_sc_hd__nor2_1 _22328_ (.A(_04923_),
    .B(_09102_),
    .Y(_01873_));
 sky130_fd_sc_hd__nor2_1 _22329_ (.A(_04932_),
    .B(_09102_),
    .Y(_01874_));
 sky130_fd_sc_hd__nor2_1 _22330_ (.A(net1142),
    .B(_09102_),
    .Y(_01875_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_712 ();
 sky130_fd_sc_hd__nor2_1 _22332_ (.A(_04951_),
    .B(_09102_),
    .Y(_01876_));
 sky130_fd_sc_hd__nor2_1 _22333_ (.A(_04794_),
    .B(_09102_),
    .Y(_01877_));
 sky130_fd_sc_hd__nor2_1 _22334_ (.A(_04960_),
    .B(_09102_),
    .Y(_01878_));
 sky130_fd_sc_hd__nor2_1 _22335_ (.A(_04974_),
    .B(_09102_),
    .Y(_01879_));
 sky130_fd_sc_hd__nor2_1 _22336_ (.A(net1137),
    .B(_09102_),
    .Y(_01880_));
 sky130_fd_sc_hd__nor2_1 _22337_ (.A(_04990_),
    .B(_09102_),
    .Y(_01881_));
 sky130_fd_sc_hd__nor2_1 _22338_ (.A(net1128),
    .B(_09102_),
    .Y(_01882_));
 sky130_fd_sc_hd__nor2_1 _22339_ (.A(_05011_),
    .B(_09102_),
    .Y(_01883_));
 sky130_fd_sc_hd__nor2_1 _22340_ (.A(_05020_),
    .B(_09102_),
    .Y(_01884_));
 sky130_fd_sc_hd__nor2_1 _22341_ (.A(_05029_),
    .B(_09102_),
    .Y(_01885_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_711 ();
 sky130_fd_sc_hd__nor2_1 _22343_ (.A(net1135),
    .B(_09102_),
    .Y(_01886_));
 sky130_fd_sc_hd__nor2_1 _22344_ (.A(_05044_),
    .B(_09102_),
    .Y(_01887_));
 sky130_fd_sc_hd__nor2_1 _22345_ (.A(_04801_),
    .B(_09102_),
    .Y(_01888_));
 sky130_fd_sc_hd__nor2_1 _22346_ (.A(_05060_),
    .B(_09102_),
    .Y(_01889_));
 sky130_fd_sc_hd__nor2_1 _22347_ (.A(_08895_),
    .B(_09102_),
    .Y(_01890_));
 sky130_fd_sc_hd__nor2_1 _22348_ (.A(_04808_),
    .B(_09102_),
    .Y(_01891_));
 sky130_fd_sc_hd__nor2_1 _22349_ (.A(_04817_),
    .B(_09102_),
    .Y(_01892_));
 sky130_fd_sc_hd__nor2_1 _22350_ (.A(_04826_),
    .B(_09102_),
    .Y(_01893_));
 sky130_fd_sc_hd__nor2_1 _22351_ (.A(_04834_),
    .B(_09102_),
    .Y(_01894_));
 sky130_fd_sc_hd__nor2_1 _22352_ (.A(_04843_),
    .B(_09102_),
    .Y(_01895_));
 sky130_fd_sc_hd__nor2_1 _22353_ (.A(_04852_),
    .B(_09102_),
    .Y(_01896_));
 sky130_fd_sc_hd__nor2_1 _22354_ (.A(_04860_),
    .B(_09102_),
    .Y(_01897_));
 sky130_fd_sc_hd__nand2_8 _22355_ (.A(_09818_),
    .B(_05474_),
    .Y(_09106_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_710 ();
 sky130_fd_sc_hd__nor2_1 _22357_ (.A(_05118_),
    .B(_09106_),
    .Y(_01898_));
 sky130_fd_sc_hd__nor2_1 _22358_ (.A(_05192_),
    .B(_09106_),
    .Y(_01899_));
 sky130_fd_sc_hd__nor2_1 _22359_ (.A(_05204_),
    .B(_09106_),
    .Y(_01900_));
 sky130_fd_sc_hd__nor2_1 _22360_ (.A(_05214_),
    .B(_09106_),
    .Y(_01901_));
 sky130_fd_sc_hd__nor2_1 _22361_ (.A(_05221_),
    .B(_09106_),
    .Y(_01902_));
 sky130_fd_sc_hd__nor2_1 _22362_ (.A(net1138),
    .B(_09106_),
    .Y(_01903_));
 sky130_fd_sc_hd__nor2_1 _22363_ (.A(_05238_),
    .B(_09106_),
    .Y(_01904_));
 sky130_fd_sc_hd__nor2_1 _22364_ (.A(_05247_),
    .B(_09106_),
    .Y(_01905_));
 sky130_fd_sc_hd__nor2_1 _22365_ (.A(_05258_),
    .B(_09106_),
    .Y(_01906_));
 sky130_fd_sc_hd__nor2_1 _22366_ (.A(net1136),
    .B(_09106_),
    .Y(_01907_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_709 ();
 sky130_fd_sc_hd__nor2_1 _22368_ (.A(_05280_),
    .B(_09106_),
    .Y(_01908_));
 sky130_fd_sc_hd__nor2_1 _22369_ (.A(_05122_),
    .B(_09106_),
    .Y(_01909_));
 sky130_fd_sc_hd__nor2_1 _22370_ (.A(_05291_),
    .B(_09106_),
    .Y(_01910_));
 sky130_fd_sc_hd__nor2_1 _22371_ (.A(_05301_),
    .B(_09106_),
    .Y(_01911_));
 sky130_fd_sc_hd__nor2_1 _22372_ (.A(_05309_),
    .B(_09106_),
    .Y(_01912_));
 sky130_fd_sc_hd__nor2_1 _22373_ (.A(_05320_),
    .B(_09106_),
    .Y(_01913_));
 sky130_fd_sc_hd__nor2_1 _22374_ (.A(net1112),
    .B(_09106_),
    .Y(_01914_));
 sky130_fd_sc_hd__nor2_1 _22375_ (.A(_05339_),
    .B(_09106_),
    .Y(_01915_));
 sky130_fd_sc_hd__nor2_1 _22376_ (.A(net1144),
    .B(_09106_),
    .Y(_01916_));
 sky130_fd_sc_hd__nor2_1 _22377_ (.A(_05358_),
    .B(_09106_),
    .Y(_01917_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_708 ();
 sky130_fd_sc_hd__nor2_1 _22379_ (.A(net1141),
    .B(_09106_),
    .Y(_01918_));
 sky130_fd_sc_hd__nor2_1 _22380_ (.A(_05380_),
    .B(_09106_),
    .Y(_01919_));
 sky130_fd_sc_hd__nor2_1 _22381_ (.A(_05126_),
    .B(_09106_),
    .Y(_01920_));
 sky130_fd_sc_hd__nor2_1 _22382_ (.A(net1114),
    .B(_09106_),
    .Y(_01921_));
 sky130_fd_sc_hd__nor2_1 _22383_ (.A(_05430_),
    .B(_09106_),
    .Y(_01922_));
 sky130_fd_sc_hd__nor2_1 _22384_ (.A(_05132_),
    .B(_09106_),
    .Y(_01923_));
 sky130_fd_sc_hd__nor2_1 _22385_ (.A(_05140_),
    .B(_09106_),
    .Y(_01924_));
 sky130_fd_sc_hd__nor2_1 _22386_ (.A(_05149_),
    .B(_09106_),
    .Y(_01925_));
 sky130_fd_sc_hd__nor2_1 _22387_ (.A(_05157_),
    .B(_09106_),
    .Y(_01926_));
 sky130_fd_sc_hd__nor2_1 _22388_ (.A(_05166_),
    .B(_09106_),
    .Y(_01927_));
 sky130_fd_sc_hd__nor2_1 _22389_ (.A(_05173_),
    .B(_09106_),
    .Y(_01928_));
 sky130_fd_sc_hd__nor2_1 _22390_ (.A(_05183_),
    .B(_09106_),
    .Y(_01929_));
 sky130_fd_sc_hd__nand2_8 _22391_ (.A(_09764_),
    .B(_05516_),
    .Y(_09110_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_707 ();
 sky130_fd_sc_hd__nor2_1 _22393_ (.A(_04790_),
    .B(_09110_),
    .Y(_01930_));
 sky130_fd_sc_hd__nor2_1 _22394_ (.A(_04871_),
    .B(_09110_),
    .Y(_01931_));
 sky130_fd_sc_hd__nor2_1 _22395_ (.A(_04883_),
    .B(_09110_),
    .Y(_01932_));
 sky130_fd_sc_hd__nor2_1 _22396_ (.A(_04892_),
    .B(_09110_),
    .Y(_01933_));
 sky130_fd_sc_hd__nor2_1 _22397_ (.A(_04899_),
    .B(_09110_),
    .Y(_01934_));
 sky130_fd_sc_hd__nor2_1 _22398_ (.A(_04906_),
    .B(_09110_),
    .Y(_01935_));
 sky130_fd_sc_hd__nor2_1 _22399_ (.A(_04913_),
    .B(_09110_),
    .Y(_01936_));
 sky130_fd_sc_hd__nor2_1 _22400_ (.A(_04923_),
    .B(_09110_),
    .Y(_01937_));
 sky130_fd_sc_hd__nor2_1 _22401_ (.A(_04932_),
    .B(_09110_),
    .Y(_01938_));
 sky130_fd_sc_hd__nor2_1 _22402_ (.A(net1142),
    .B(_09110_),
    .Y(_01939_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_706 ();
 sky130_fd_sc_hd__nor2_1 _22404_ (.A(_04951_),
    .B(_09110_),
    .Y(_01940_));
 sky130_fd_sc_hd__nor2_1 _22405_ (.A(_04794_),
    .B(_09110_),
    .Y(_01941_));
 sky130_fd_sc_hd__nor2_1 _22406_ (.A(_04960_),
    .B(_09110_),
    .Y(_01942_));
 sky130_fd_sc_hd__nor2_1 _22407_ (.A(_04974_),
    .B(_09110_),
    .Y(_01943_));
 sky130_fd_sc_hd__nor2_1 _22408_ (.A(_04984_),
    .B(_09110_),
    .Y(_01944_));
 sky130_fd_sc_hd__nor2_1 _22409_ (.A(_04990_),
    .B(_09110_),
    .Y(_01945_));
 sky130_fd_sc_hd__nor2_1 _22410_ (.A(net1128),
    .B(_09110_),
    .Y(_01946_));
 sky130_fd_sc_hd__nor2_1 _22411_ (.A(_05011_),
    .B(_09110_),
    .Y(_01947_));
 sky130_fd_sc_hd__nor2_1 _22412_ (.A(_05020_),
    .B(_09110_),
    .Y(_01948_));
 sky130_fd_sc_hd__nor2_1 _22413_ (.A(_05029_),
    .B(_09110_),
    .Y(_01949_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_705 ();
 sky130_fd_sc_hd__nor2_1 _22415_ (.A(_05035_),
    .B(_09110_),
    .Y(_01950_));
 sky130_fd_sc_hd__nor2_1 _22416_ (.A(_05044_),
    .B(_09110_),
    .Y(_01951_));
 sky130_fd_sc_hd__nor2_1 _22417_ (.A(_04801_),
    .B(_09110_),
    .Y(_01952_));
 sky130_fd_sc_hd__nor2_1 _22418_ (.A(_05060_),
    .B(_09110_),
    .Y(_01953_));
 sky130_fd_sc_hd__nor2_1 _22419_ (.A(_08895_),
    .B(_09110_),
    .Y(_01954_));
 sky130_fd_sc_hd__nor2_1 _22420_ (.A(_04808_),
    .B(_09110_),
    .Y(_01955_));
 sky130_fd_sc_hd__nor2_1 _22421_ (.A(_04817_),
    .B(_09110_),
    .Y(_01956_));
 sky130_fd_sc_hd__nor2_1 _22422_ (.A(_04826_),
    .B(_09110_),
    .Y(_01957_));
 sky130_fd_sc_hd__nor2_1 _22423_ (.A(_04834_),
    .B(_09110_),
    .Y(_01958_));
 sky130_fd_sc_hd__nor2_1 _22424_ (.A(_04843_),
    .B(_09110_),
    .Y(_01959_));
 sky130_fd_sc_hd__nor2_1 _22425_ (.A(_04852_),
    .B(_09110_),
    .Y(_01960_));
 sky130_fd_sc_hd__nor2_1 _22426_ (.A(_04860_),
    .B(_09110_),
    .Y(_01961_));
 sky130_fd_sc_hd__nand2_8 _22427_ (.A(_09818_),
    .B(_05557_),
    .Y(_09114_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_704 ();
 sky130_fd_sc_hd__nor2_1 _22429_ (.A(_05118_),
    .B(_09114_),
    .Y(_01962_));
 sky130_fd_sc_hd__nor2_1 _22430_ (.A(_05192_),
    .B(_09114_),
    .Y(_01963_));
 sky130_fd_sc_hd__nor2_1 _22431_ (.A(_05204_),
    .B(_09114_),
    .Y(_01964_));
 sky130_fd_sc_hd__nor2_1 _22432_ (.A(_05214_),
    .B(_09114_),
    .Y(_01965_));
 sky130_fd_sc_hd__nor2_1 _22433_ (.A(_05221_),
    .B(_09114_),
    .Y(_01966_));
 sky130_fd_sc_hd__nor2_1 _22434_ (.A(net1138),
    .B(_09114_),
    .Y(_01967_));
 sky130_fd_sc_hd__nor2_1 _22435_ (.A(_05238_),
    .B(_09114_),
    .Y(_01968_));
 sky130_fd_sc_hd__nor2_1 _22436_ (.A(net1140),
    .B(_09114_),
    .Y(_01969_));
 sky130_fd_sc_hd__nor2_1 _22437_ (.A(_05258_),
    .B(_09114_),
    .Y(_01970_));
 sky130_fd_sc_hd__nor2_1 _22438_ (.A(net1136),
    .B(_09114_),
    .Y(_01971_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_703 ();
 sky130_fd_sc_hd__nor2_1 _22440_ (.A(_05280_),
    .B(_09114_),
    .Y(_01972_));
 sky130_fd_sc_hd__nor2_1 _22441_ (.A(_05122_),
    .B(_09114_),
    .Y(_01973_));
 sky130_fd_sc_hd__nor2_1 _22442_ (.A(_05291_),
    .B(_09114_),
    .Y(_01974_));
 sky130_fd_sc_hd__nor2_1 _22443_ (.A(_05301_),
    .B(_09114_),
    .Y(_01975_));
 sky130_fd_sc_hd__nor2_1 _22444_ (.A(_05309_),
    .B(_09114_),
    .Y(_01976_));
 sky130_fd_sc_hd__nor2_1 _22445_ (.A(_05320_),
    .B(_09114_),
    .Y(_01977_));
 sky130_fd_sc_hd__nor2_1 _22446_ (.A(net1112),
    .B(_09114_),
    .Y(_01978_));
 sky130_fd_sc_hd__nor2_1 _22447_ (.A(_05339_),
    .B(_09114_),
    .Y(_01979_));
 sky130_fd_sc_hd__nor2_1 _22448_ (.A(net1144),
    .B(_09114_),
    .Y(_01980_));
 sky130_fd_sc_hd__nor2_1 _22449_ (.A(_05358_),
    .B(_09114_),
    .Y(_01981_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_702 ();
 sky130_fd_sc_hd__nor2_1 _22451_ (.A(net1113),
    .B(_09114_),
    .Y(_01982_));
 sky130_fd_sc_hd__nor2_1 _22452_ (.A(_05380_),
    .B(_09114_),
    .Y(_01983_));
 sky130_fd_sc_hd__nor2_1 _22453_ (.A(_05126_),
    .B(_09114_),
    .Y(_01984_));
 sky130_fd_sc_hd__nor2_1 _22454_ (.A(net1143),
    .B(_09114_),
    .Y(_01985_));
 sky130_fd_sc_hd__nor2_1 _22455_ (.A(_05430_),
    .B(_09114_),
    .Y(_01986_));
 sky130_fd_sc_hd__nor2_1 _22456_ (.A(_05132_),
    .B(_09114_),
    .Y(_01987_));
 sky130_fd_sc_hd__nor2_1 _22457_ (.A(_05140_),
    .B(_09114_),
    .Y(_01988_));
 sky130_fd_sc_hd__nor2_1 _22458_ (.A(_05149_),
    .B(_09114_),
    .Y(_01989_));
 sky130_fd_sc_hd__nor2_1 _22459_ (.A(_05157_),
    .B(_09114_),
    .Y(_01990_));
 sky130_fd_sc_hd__nor2_1 _22460_ (.A(_05166_),
    .B(_09114_),
    .Y(_01991_));
 sky130_fd_sc_hd__nor2_1 _22461_ (.A(_05173_),
    .B(_09114_),
    .Y(_01992_));
 sky130_fd_sc_hd__nor2_1 _22462_ (.A(_05183_),
    .B(_09114_),
    .Y(_01993_));
 sky130_fd_sc_hd__nand2_8 _22463_ (.A(_09764_),
    .B(_05598_),
    .Y(_09118_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_701 ();
 sky130_fd_sc_hd__nor2_1 _22465_ (.A(_04790_),
    .B(_09118_),
    .Y(_01994_));
 sky130_fd_sc_hd__nor2_1 _22466_ (.A(_04871_),
    .B(_09118_),
    .Y(_01995_));
 sky130_fd_sc_hd__nor2_1 _22467_ (.A(_04883_),
    .B(_09118_),
    .Y(_01996_));
 sky130_fd_sc_hd__nor2_1 _22468_ (.A(_04892_),
    .B(_09118_),
    .Y(_01997_));
 sky130_fd_sc_hd__nor2_1 _22469_ (.A(_04899_),
    .B(_09118_),
    .Y(_01998_));
 sky130_fd_sc_hd__nor2_1 _22470_ (.A(_04906_),
    .B(_09118_),
    .Y(_01999_));
 sky130_fd_sc_hd__nor2_1 _22471_ (.A(_04913_),
    .B(_09118_),
    .Y(_02000_));
 sky130_fd_sc_hd__nor2_1 _22472_ (.A(_04923_),
    .B(_09118_),
    .Y(_02001_));
 sky130_fd_sc_hd__nor2_1 _22473_ (.A(_04932_),
    .B(_09118_),
    .Y(_02002_));
 sky130_fd_sc_hd__nor2_1 _22474_ (.A(net1142),
    .B(_09118_),
    .Y(_02003_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_700 ();
 sky130_fd_sc_hd__nor2_1 _22476_ (.A(_04951_),
    .B(_09118_),
    .Y(_02004_));
 sky130_fd_sc_hd__nor2_1 _22477_ (.A(_04794_),
    .B(_09118_),
    .Y(_02005_));
 sky130_fd_sc_hd__nor2_1 _22478_ (.A(_04960_),
    .B(_09118_),
    .Y(_02006_));
 sky130_fd_sc_hd__nor2_1 _22479_ (.A(_04974_),
    .B(_09118_),
    .Y(_02007_));
 sky130_fd_sc_hd__nor2_1 _22480_ (.A(net1137),
    .B(_09118_),
    .Y(_02008_));
 sky130_fd_sc_hd__nor2_1 _22481_ (.A(_04990_),
    .B(_09118_),
    .Y(_02009_));
 sky130_fd_sc_hd__nor2_1 _22482_ (.A(net1128),
    .B(_09118_),
    .Y(_02010_));
 sky130_fd_sc_hd__nor2_1 _22483_ (.A(_05011_),
    .B(_09118_),
    .Y(_02011_));
 sky130_fd_sc_hd__nor2_1 _22484_ (.A(net1139),
    .B(_09118_),
    .Y(_02012_));
 sky130_fd_sc_hd__nor2_1 _22485_ (.A(_05029_),
    .B(_09118_),
    .Y(_02013_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_699 ();
 sky130_fd_sc_hd__nor2_1 _22487_ (.A(net1135),
    .B(_09118_),
    .Y(_02014_));
 sky130_fd_sc_hd__nor2_1 _22488_ (.A(_05044_),
    .B(_09118_),
    .Y(_02015_));
 sky130_fd_sc_hd__nor2_1 _22489_ (.A(_04801_),
    .B(_09118_),
    .Y(_02016_));
 sky130_fd_sc_hd__nor2_1 _22490_ (.A(_05060_),
    .B(_09118_),
    .Y(_02017_));
 sky130_fd_sc_hd__nor2_1 _22491_ (.A(_08895_),
    .B(_09118_),
    .Y(_02018_));
 sky130_fd_sc_hd__nor2_1 _22492_ (.A(_04808_),
    .B(_09118_),
    .Y(_02019_));
 sky130_fd_sc_hd__nor2_1 _22493_ (.A(_04817_),
    .B(_09118_),
    .Y(_02020_));
 sky130_fd_sc_hd__nor2_1 _22494_ (.A(_04826_),
    .B(_09118_),
    .Y(_02021_));
 sky130_fd_sc_hd__nor2_1 _22495_ (.A(_04834_),
    .B(_09118_),
    .Y(_02022_));
 sky130_fd_sc_hd__nor2_1 _22496_ (.A(_04843_),
    .B(_09118_),
    .Y(_02023_));
 sky130_fd_sc_hd__nor2_1 _22497_ (.A(_04852_),
    .B(_09118_),
    .Y(_02024_));
 sky130_fd_sc_hd__nor2_1 _22498_ (.A(_04860_),
    .B(_09118_),
    .Y(_02025_));
 sky130_fd_sc_hd__nand2_8 _22499_ (.A(_09818_),
    .B(_05951_),
    .Y(_09122_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_698 ();
 sky130_fd_sc_hd__nor2_1 _22501_ (.A(_05118_),
    .B(_09122_),
    .Y(_02026_));
 sky130_fd_sc_hd__nor2_1 _22502_ (.A(_05192_),
    .B(_09122_),
    .Y(_02027_));
 sky130_fd_sc_hd__nor2_1 _22503_ (.A(_05204_),
    .B(_09122_),
    .Y(_02028_));
 sky130_fd_sc_hd__nor2_1 _22504_ (.A(_05214_),
    .B(_09122_),
    .Y(_02029_));
 sky130_fd_sc_hd__nor2_1 _22505_ (.A(_05221_),
    .B(_09122_),
    .Y(_02030_));
 sky130_fd_sc_hd__nor2_1 _22506_ (.A(_05228_),
    .B(_09122_),
    .Y(_02031_));
 sky130_fd_sc_hd__nor2_1 _22507_ (.A(_05238_),
    .B(_09122_),
    .Y(_02032_));
 sky130_fd_sc_hd__nor2_1 _22508_ (.A(_05247_),
    .B(_09122_),
    .Y(_02033_));
 sky130_fd_sc_hd__nor2_1 _22509_ (.A(_05258_),
    .B(_09122_),
    .Y(_02034_));
 sky130_fd_sc_hd__nor2_1 _22510_ (.A(net1136),
    .B(_09122_),
    .Y(_02035_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_697 ();
 sky130_fd_sc_hd__nor2_1 _22512_ (.A(_05280_),
    .B(_09122_),
    .Y(_02036_));
 sky130_fd_sc_hd__nor2_1 _22513_ (.A(_05122_),
    .B(_09122_),
    .Y(_02037_));
 sky130_fd_sc_hd__nor2_1 _22514_ (.A(_05291_),
    .B(_09122_),
    .Y(_02038_));
 sky130_fd_sc_hd__nor2_1 _22515_ (.A(_05301_),
    .B(_09122_),
    .Y(_02039_));
 sky130_fd_sc_hd__nor2_1 _22516_ (.A(_05309_),
    .B(_09122_),
    .Y(_02040_));
 sky130_fd_sc_hd__nor2_1 _22517_ (.A(_05320_),
    .B(_09122_),
    .Y(_02041_));
 sky130_fd_sc_hd__nor2_1 _22518_ (.A(net1112),
    .B(_09122_),
    .Y(_02042_));
 sky130_fd_sc_hd__nor2_1 _22519_ (.A(_05339_),
    .B(_09122_),
    .Y(_02043_));
 sky130_fd_sc_hd__nor2_1 _22520_ (.A(_05347_),
    .B(_09122_),
    .Y(_02044_));
 sky130_fd_sc_hd__nor2_1 _22521_ (.A(_05358_),
    .B(_09122_),
    .Y(_02045_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_696 ();
 sky130_fd_sc_hd__nor2_1 _22523_ (.A(net1134),
    .B(_09122_),
    .Y(_02046_));
 sky130_fd_sc_hd__nor2_1 _22524_ (.A(_05380_),
    .B(_09122_),
    .Y(_02047_));
 sky130_fd_sc_hd__nor2_1 _22525_ (.A(_05126_),
    .B(_09122_),
    .Y(_02048_));
 sky130_fd_sc_hd__nor2_1 _22526_ (.A(net1114),
    .B(_09122_),
    .Y(_02049_));
 sky130_fd_sc_hd__nor2_1 _22527_ (.A(_05430_),
    .B(_09122_),
    .Y(_02050_));
 sky130_fd_sc_hd__nor2_1 _22528_ (.A(_05132_),
    .B(_09122_),
    .Y(_02051_));
 sky130_fd_sc_hd__nor2_1 _22529_ (.A(_05140_),
    .B(_09122_),
    .Y(_02052_));
 sky130_fd_sc_hd__nor2_1 _22530_ (.A(_05149_),
    .B(_09122_),
    .Y(_02053_));
 sky130_fd_sc_hd__nor2_1 _22531_ (.A(_05157_),
    .B(_09122_),
    .Y(_02054_));
 sky130_fd_sc_hd__nor2_1 _22532_ (.A(_05166_),
    .B(_09122_),
    .Y(_02055_));
 sky130_fd_sc_hd__nor2_1 _22533_ (.A(_05173_),
    .B(_09122_),
    .Y(_02056_));
 sky130_fd_sc_hd__nor2_1 _22534_ (.A(_05183_),
    .B(_09122_),
    .Y(_02057_));
 sky130_fd_sc_hd__nand2_8 _22535_ (.A(_09771_),
    .B(_04784_),
    .Y(_09126_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_695 ();
 sky130_fd_sc_hd__nor2_1 _22537_ (.A(_04790_),
    .B(_09126_),
    .Y(_02058_));
 sky130_fd_sc_hd__nor2_1 _22538_ (.A(_04871_),
    .B(_09126_),
    .Y(_02059_));
 sky130_fd_sc_hd__nor2_1 _22539_ (.A(_04883_),
    .B(_09126_),
    .Y(_02060_));
 sky130_fd_sc_hd__nor2_1 _22540_ (.A(_04892_),
    .B(_09126_),
    .Y(_02061_));
 sky130_fd_sc_hd__nor2_1 _22541_ (.A(_04899_),
    .B(_09126_),
    .Y(_02062_));
 sky130_fd_sc_hd__nor2_1 _22542_ (.A(_04906_),
    .B(_09126_),
    .Y(_02063_));
 sky130_fd_sc_hd__nor2_1 _22543_ (.A(_04913_),
    .B(_09126_),
    .Y(_02064_));
 sky130_fd_sc_hd__nor2_1 _22544_ (.A(_04923_),
    .B(_09126_),
    .Y(_02065_));
 sky130_fd_sc_hd__nor2_1 _22545_ (.A(_04932_),
    .B(_09126_),
    .Y(_02066_));
 sky130_fd_sc_hd__nor2_1 _22546_ (.A(net1142),
    .B(_09126_),
    .Y(_02067_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_694 ();
 sky130_fd_sc_hd__nor2_1 _22548_ (.A(_04951_),
    .B(_09126_),
    .Y(_02068_));
 sky130_fd_sc_hd__nor2_1 _22549_ (.A(_04794_),
    .B(_09126_),
    .Y(_02069_));
 sky130_fd_sc_hd__nor2_1 _22550_ (.A(_04960_),
    .B(_09126_),
    .Y(_02070_));
 sky130_fd_sc_hd__nor2_1 _22551_ (.A(_04974_),
    .B(_09126_),
    .Y(_02071_));
 sky130_fd_sc_hd__nor2_1 _22552_ (.A(net1137),
    .B(_09126_),
    .Y(_02072_));
 sky130_fd_sc_hd__nor2_1 _22553_ (.A(_04990_),
    .B(_09126_),
    .Y(_02073_));
 sky130_fd_sc_hd__nor2_1 _22554_ (.A(net1128),
    .B(_09126_),
    .Y(_02074_));
 sky130_fd_sc_hd__nor2_1 _22555_ (.A(_05011_),
    .B(_09126_),
    .Y(_02075_));
 sky130_fd_sc_hd__nor2_1 _22556_ (.A(_05020_),
    .B(_09126_),
    .Y(_02076_));
 sky130_fd_sc_hd__nor2_1 _22557_ (.A(_05029_),
    .B(_09126_),
    .Y(_02077_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_693 ();
 sky130_fd_sc_hd__nor2_1 _22559_ (.A(_05035_),
    .B(_09126_),
    .Y(_02078_));
 sky130_fd_sc_hd__nor2_1 _22560_ (.A(_05044_),
    .B(_09126_),
    .Y(_02079_));
 sky130_fd_sc_hd__nor2_1 _22561_ (.A(_04801_),
    .B(_09126_),
    .Y(_02080_));
 sky130_fd_sc_hd__nor2_1 _22562_ (.A(_05060_),
    .B(_09126_),
    .Y(_02081_));
 sky130_fd_sc_hd__nor2_1 _22563_ (.A(_08895_),
    .B(_09126_),
    .Y(_02082_));
 sky130_fd_sc_hd__nor2_1 _22564_ (.A(_04808_),
    .B(_09126_),
    .Y(_02083_));
 sky130_fd_sc_hd__nor2_1 _22565_ (.A(_04817_),
    .B(_09126_),
    .Y(_02084_));
 sky130_fd_sc_hd__nor2_1 _22566_ (.A(_04826_),
    .B(_09126_),
    .Y(_02085_));
 sky130_fd_sc_hd__nor2_1 _22567_ (.A(_04834_),
    .B(_09126_),
    .Y(_02086_));
 sky130_fd_sc_hd__nor2_1 _22568_ (.A(_04843_),
    .B(_09126_),
    .Y(_02087_));
 sky130_fd_sc_hd__nor2_1 _22569_ (.A(_04852_),
    .B(_09126_),
    .Y(_02088_));
 sky130_fd_sc_hd__nor2_1 _22570_ (.A(_04860_),
    .B(_09126_),
    .Y(_02089_));
 sky130_fd_sc_hd__nand2_8 _22571_ (.A(_09825_),
    .B(_05115_),
    .Y(_09130_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_692 ();
 sky130_fd_sc_hd__nor2_1 _22573_ (.A(_05118_),
    .B(_09130_),
    .Y(_02090_));
 sky130_fd_sc_hd__nor2_1 _22574_ (.A(_05192_),
    .B(_09130_),
    .Y(_02091_));
 sky130_fd_sc_hd__nor2_1 _22575_ (.A(_05204_),
    .B(_09130_),
    .Y(_02092_));
 sky130_fd_sc_hd__nor2_1 _22576_ (.A(_05214_),
    .B(_09130_),
    .Y(_02093_));
 sky130_fd_sc_hd__nor2_1 _22577_ (.A(_05221_),
    .B(_09130_),
    .Y(_02094_));
 sky130_fd_sc_hd__nor2_1 _22578_ (.A(_05228_),
    .B(_09130_),
    .Y(_02095_));
 sky130_fd_sc_hd__nor2_1 _22579_ (.A(_05238_),
    .B(_09130_),
    .Y(_02096_));
 sky130_fd_sc_hd__nor2_1 _22580_ (.A(net1140),
    .B(_09130_),
    .Y(_02097_));
 sky130_fd_sc_hd__nor2_1 _22581_ (.A(_05258_),
    .B(_09130_),
    .Y(_02098_));
 sky130_fd_sc_hd__nor2_1 _22582_ (.A(net1136),
    .B(_09130_),
    .Y(_02099_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_691 ();
 sky130_fd_sc_hd__nor2_1 _22584_ (.A(_05280_),
    .B(_09130_),
    .Y(_02100_));
 sky130_fd_sc_hd__nor2_1 _22585_ (.A(_05122_),
    .B(_09130_),
    .Y(_02101_));
 sky130_fd_sc_hd__nor2_1 _22586_ (.A(_05291_),
    .B(_09130_),
    .Y(_02102_));
 sky130_fd_sc_hd__nor2_1 _22587_ (.A(_05301_),
    .B(_09130_),
    .Y(_02103_));
 sky130_fd_sc_hd__nor2_1 _22588_ (.A(_05309_),
    .B(_09130_),
    .Y(_02104_));
 sky130_fd_sc_hd__nor2_1 _22589_ (.A(_05320_),
    .B(_09130_),
    .Y(_02105_));
 sky130_fd_sc_hd__nor2_1 _22590_ (.A(net1112),
    .B(_09130_),
    .Y(_02106_));
 sky130_fd_sc_hd__nor2_1 _22591_ (.A(_05339_),
    .B(_09130_),
    .Y(_02107_));
 sky130_fd_sc_hd__nor2_1 _22592_ (.A(net1144),
    .B(_09130_),
    .Y(_02108_));
 sky130_fd_sc_hd__nor2_1 _22593_ (.A(_05358_),
    .B(_09130_),
    .Y(_02109_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_690 ();
 sky130_fd_sc_hd__nor2_1 _22595_ (.A(net1113),
    .B(_09130_),
    .Y(_02110_));
 sky130_fd_sc_hd__nor2_1 _22596_ (.A(_05380_),
    .B(_09130_),
    .Y(_02111_));
 sky130_fd_sc_hd__nor2_1 _22597_ (.A(_05126_),
    .B(_09130_),
    .Y(_02112_));
 sky130_fd_sc_hd__nor2_1 _22598_ (.A(net1114),
    .B(_09130_),
    .Y(_02113_));
 sky130_fd_sc_hd__nor2_1 _22599_ (.A(_05430_),
    .B(_09130_),
    .Y(_02114_));
 sky130_fd_sc_hd__nor2_1 _22600_ (.A(_05132_),
    .B(_09130_),
    .Y(_02115_));
 sky130_fd_sc_hd__nor2_1 _22601_ (.A(_05140_),
    .B(_09130_),
    .Y(_02116_));
 sky130_fd_sc_hd__nor2_1 _22602_ (.A(_05149_),
    .B(_09130_),
    .Y(_02117_));
 sky130_fd_sc_hd__nor2_1 _22603_ (.A(_05157_),
    .B(_09130_),
    .Y(_02118_));
 sky130_fd_sc_hd__nor2_1 _22604_ (.A(_05166_),
    .B(_09130_),
    .Y(_02119_));
 sky130_fd_sc_hd__nor2_1 _22605_ (.A(_05173_),
    .B(_09130_),
    .Y(_02120_));
 sky130_fd_sc_hd__nor2_1 _22606_ (.A(_05183_),
    .B(_09130_),
    .Y(_02121_));
 sky130_fd_sc_hd__nand2_8 _22607_ (.A(_09771_),
    .B(_05433_),
    .Y(_09134_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_689 ();
 sky130_fd_sc_hd__nor2_1 _22609_ (.A(_04790_),
    .B(_09134_),
    .Y(_02122_));
 sky130_fd_sc_hd__nor2_1 _22610_ (.A(_04871_),
    .B(_09134_),
    .Y(_02123_));
 sky130_fd_sc_hd__nor2_1 _22611_ (.A(_04883_),
    .B(_09134_),
    .Y(_02124_));
 sky130_fd_sc_hd__nor2_1 _22612_ (.A(_04892_),
    .B(_09134_),
    .Y(_02125_));
 sky130_fd_sc_hd__nor2_1 _22613_ (.A(_04899_),
    .B(_09134_),
    .Y(_02126_));
 sky130_fd_sc_hd__nor2_1 _22614_ (.A(_04906_),
    .B(_09134_),
    .Y(_02127_));
 sky130_fd_sc_hd__nor2_1 _22615_ (.A(_04913_),
    .B(_09134_),
    .Y(_02128_));
 sky130_fd_sc_hd__nor2_1 _22616_ (.A(_04923_),
    .B(_09134_),
    .Y(_02129_));
 sky130_fd_sc_hd__nor2_1 _22617_ (.A(_04932_),
    .B(_09134_),
    .Y(_02130_));
 sky130_fd_sc_hd__nor2_1 _22618_ (.A(net1142),
    .B(_09134_),
    .Y(_02131_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_688 ();
 sky130_fd_sc_hd__nor2_1 _22620_ (.A(_04951_),
    .B(_09134_),
    .Y(_02132_));
 sky130_fd_sc_hd__nor2_1 _22621_ (.A(_04794_),
    .B(_09134_),
    .Y(_02133_));
 sky130_fd_sc_hd__nor2_1 _22622_ (.A(_04960_),
    .B(_09134_),
    .Y(_02134_));
 sky130_fd_sc_hd__nor2_1 _22623_ (.A(_04974_),
    .B(_09134_),
    .Y(_02135_));
 sky130_fd_sc_hd__nor2_1 _22624_ (.A(net1137),
    .B(_09134_),
    .Y(_02136_));
 sky130_fd_sc_hd__nor2_1 _22625_ (.A(_04990_),
    .B(_09134_),
    .Y(_02137_));
 sky130_fd_sc_hd__nor2_1 _22626_ (.A(net1128),
    .B(_09134_),
    .Y(_02138_));
 sky130_fd_sc_hd__nor2_1 _22627_ (.A(_05011_),
    .B(_09134_),
    .Y(_02139_));
 sky130_fd_sc_hd__nor2_1 _22628_ (.A(net1139),
    .B(_09134_),
    .Y(_02140_));
 sky130_fd_sc_hd__nor2_1 _22629_ (.A(_05029_),
    .B(_09134_),
    .Y(_02141_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_687 ();
 sky130_fd_sc_hd__nor2_1 _22631_ (.A(net1135),
    .B(_09134_),
    .Y(_02142_));
 sky130_fd_sc_hd__nor2_1 _22632_ (.A(_05044_),
    .B(_09134_),
    .Y(_02143_));
 sky130_fd_sc_hd__nor2_1 _22633_ (.A(_04801_),
    .B(_09134_),
    .Y(_02144_));
 sky130_fd_sc_hd__nor2_1 _22634_ (.A(_05060_),
    .B(_09134_),
    .Y(_02145_));
 sky130_fd_sc_hd__nor2_1 _22635_ (.A(_08895_),
    .B(_09134_),
    .Y(_02146_));
 sky130_fd_sc_hd__nor2_1 _22636_ (.A(_04808_),
    .B(_09134_),
    .Y(_02147_));
 sky130_fd_sc_hd__nor2_1 _22637_ (.A(_04817_),
    .B(_09134_),
    .Y(_02148_));
 sky130_fd_sc_hd__nor2_1 _22638_ (.A(_04826_),
    .B(_09134_),
    .Y(_02149_));
 sky130_fd_sc_hd__nor2_1 _22639_ (.A(_04834_),
    .B(_09134_),
    .Y(_02150_));
 sky130_fd_sc_hd__nor2_1 _22640_ (.A(_04843_),
    .B(_09134_),
    .Y(_02151_));
 sky130_fd_sc_hd__nor2_1 _22641_ (.A(_04852_),
    .B(_09134_),
    .Y(_02152_));
 sky130_fd_sc_hd__nor2_1 _22642_ (.A(_04860_),
    .B(_09134_),
    .Y(_02153_));
 sky130_fd_sc_hd__nand2_8 _22643_ (.A(_09825_),
    .B(_05474_),
    .Y(_09138_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_686 ();
 sky130_fd_sc_hd__nor2_1 _22645_ (.A(_05118_),
    .B(_09138_),
    .Y(_02154_));
 sky130_fd_sc_hd__nor2_1 _22646_ (.A(_05192_),
    .B(_09138_),
    .Y(_02155_));
 sky130_fd_sc_hd__nor2_1 _22647_ (.A(_05204_),
    .B(_09138_),
    .Y(_02156_));
 sky130_fd_sc_hd__nor2_1 _22648_ (.A(_05214_),
    .B(_09138_),
    .Y(_02157_));
 sky130_fd_sc_hd__nor2_1 _22649_ (.A(_05221_),
    .B(_09138_),
    .Y(_02158_));
 sky130_fd_sc_hd__nor2_1 _22650_ (.A(net1138),
    .B(_09138_),
    .Y(_02159_));
 sky130_fd_sc_hd__nor2_1 _22651_ (.A(_05238_),
    .B(_09138_),
    .Y(_02160_));
 sky130_fd_sc_hd__nor2_1 _22652_ (.A(net1140),
    .B(_09138_),
    .Y(_02161_));
 sky130_fd_sc_hd__nor2_1 _22653_ (.A(_05258_),
    .B(_09138_),
    .Y(_02162_));
 sky130_fd_sc_hd__nor2_1 _22654_ (.A(_05267_),
    .B(_09138_),
    .Y(_02163_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_685 ();
 sky130_fd_sc_hd__nor2_1 _22656_ (.A(_05280_),
    .B(_09138_),
    .Y(_02164_));
 sky130_fd_sc_hd__nor2_1 _22657_ (.A(_05122_),
    .B(_09138_),
    .Y(_02165_));
 sky130_fd_sc_hd__nor2_1 _22658_ (.A(_05291_),
    .B(_09138_),
    .Y(_02166_));
 sky130_fd_sc_hd__nor2_1 _22659_ (.A(_05301_),
    .B(_09138_),
    .Y(_02167_));
 sky130_fd_sc_hd__nor2_1 _22660_ (.A(_05309_),
    .B(_09138_),
    .Y(_02168_));
 sky130_fd_sc_hd__nor2_1 _22661_ (.A(_05320_),
    .B(_09138_),
    .Y(_02169_));
 sky130_fd_sc_hd__nor2_1 _22662_ (.A(net1112),
    .B(_09138_),
    .Y(_02170_));
 sky130_fd_sc_hd__nor2_1 _22663_ (.A(_05339_),
    .B(_09138_),
    .Y(_02171_));
 sky130_fd_sc_hd__nor2_1 _22664_ (.A(net1144),
    .B(_09138_),
    .Y(_02172_));
 sky130_fd_sc_hd__nor2_1 _22665_ (.A(_05358_),
    .B(_09138_),
    .Y(_02173_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_684 ();
 sky130_fd_sc_hd__nor2_1 _22667_ (.A(net1113),
    .B(_09138_),
    .Y(_02174_));
 sky130_fd_sc_hd__nor2_1 _22668_ (.A(_05380_),
    .B(_09138_),
    .Y(_02175_));
 sky130_fd_sc_hd__nor2_1 _22669_ (.A(_05126_),
    .B(_09138_),
    .Y(_02176_));
 sky130_fd_sc_hd__nor2_1 _22670_ (.A(net1143),
    .B(_09138_),
    .Y(_02177_));
 sky130_fd_sc_hd__nor2_1 _22671_ (.A(_05430_),
    .B(_09138_),
    .Y(_02178_));
 sky130_fd_sc_hd__nor2_1 _22672_ (.A(_05132_),
    .B(_09138_),
    .Y(_02179_));
 sky130_fd_sc_hd__nor2_1 _22673_ (.A(_05140_),
    .B(_09138_),
    .Y(_02180_));
 sky130_fd_sc_hd__nor2_1 _22674_ (.A(_05149_),
    .B(_09138_),
    .Y(_02181_));
 sky130_fd_sc_hd__nor2_1 _22675_ (.A(_05157_),
    .B(_09138_),
    .Y(_02182_));
 sky130_fd_sc_hd__nor2_1 _22676_ (.A(_05166_),
    .B(_09138_),
    .Y(_02183_));
 sky130_fd_sc_hd__nor2_1 _22677_ (.A(_05173_),
    .B(_09138_),
    .Y(_02184_));
 sky130_fd_sc_hd__nor2_1 _22678_ (.A(_05183_),
    .B(_09138_),
    .Y(_02185_));
 sky130_fd_sc_hd__nand2_8 _22679_ (.A(_09771_),
    .B(_05516_),
    .Y(_09142_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_683 ();
 sky130_fd_sc_hd__nor2_1 _22681_ (.A(_04790_),
    .B(_09142_),
    .Y(_02186_));
 sky130_fd_sc_hd__nor2_1 _22682_ (.A(_04871_),
    .B(_09142_),
    .Y(_02187_));
 sky130_fd_sc_hd__nor2_1 _22683_ (.A(_04883_),
    .B(_09142_),
    .Y(_02188_));
 sky130_fd_sc_hd__nor2_1 _22684_ (.A(_04892_),
    .B(_09142_),
    .Y(_02189_));
 sky130_fd_sc_hd__nor2_1 _22685_ (.A(_04899_),
    .B(_09142_),
    .Y(_02190_));
 sky130_fd_sc_hd__nor2_1 _22686_ (.A(_04906_),
    .B(_09142_),
    .Y(_02191_));
 sky130_fd_sc_hd__nor2_1 _22687_ (.A(_04913_),
    .B(_09142_),
    .Y(_02192_));
 sky130_fd_sc_hd__nor2_1 _22688_ (.A(_04923_),
    .B(_09142_),
    .Y(_02193_));
 sky130_fd_sc_hd__nor2_1 _22689_ (.A(_04932_),
    .B(_09142_),
    .Y(_02194_));
 sky130_fd_sc_hd__nor2_1 _22690_ (.A(net1142),
    .B(_09142_),
    .Y(_02195_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_682 ();
 sky130_fd_sc_hd__nor2_1 _22692_ (.A(_04951_),
    .B(_09142_),
    .Y(_02196_));
 sky130_fd_sc_hd__nor2_1 _22693_ (.A(_04794_),
    .B(_09142_),
    .Y(_02197_));
 sky130_fd_sc_hd__nor2_1 _22694_ (.A(_04960_),
    .B(_09142_),
    .Y(_02198_));
 sky130_fd_sc_hd__nor2_1 _22695_ (.A(_04974_),
    .B(_09142_),
    .Y(_02199_));
 sky130_fd_sc_hd__nor2_1 _22696_ (.A(net1137),
    .B(_09142_),
    .Y(_02200_));
 sky130_fd_sc_hd__nor2_1 _22697_ (.A(_04990_),
    .B(_09142_),
    .Y(_02201_));
 sky130_fd_sc_hd__nor2_1 _22698_ (.A(net1128),
    .B(_09142_),
    .Y(_02202_));
 sky130_fd_sc_hd__nor2_1 _22699_ (.A(_05011_),
    .B(_09142_),
    .Y(_02203_));
 sky130_fd_sc_hd__nor2_1 _22700_ (.A(net1139),
    .B(_09142_),
    .Y(_02204_));
 sky130_fd_sc_hd__nor2_1 _22701_ (.A(_05029_),
    .B(_09142_),
    .Y(_02205_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_681 ();
 sky130_fd_sc_hd__nor2_1 _22703_ (.A(net1135),
    .B(_09142_),
    .Y(_02206_));
 sky130_fd_sc_hd__nor2_1 _22704_ (.A(_05044_),
    .B(_09142_),
    .Y(_02207_));
 sky130_fd_sc_hd__nor2_1 _22705_ (.A(_04801_),
    .B(_09142_),
    .Y(_02208_));
 sky130_fd_sc_hd__nor2_1 _22706_ (.A(_05060_),
    .B(_09142_),
    .Y(_02209_));
 sky130_fd_sc_hd__nor2_1 _22707_ (.A(_08895_),
    .B(_09142_),
    .Y(_02210_));
 sky130_fd_sc_hd__nor2_1 _22708_ (.A(_04808_),
    .B(_09142_),
    .Y(_02211_));
 sky130_fd_sc_hd__nor2_1 _22709_ (.A(_04817_),
    .B(_09142_),
    .Y(_02212_));
 sky130_fd_sc_hd__nor2_1 _22710_ (.A(_04826_),
    .B(_09142_),
    .Y(_02213_));
 sky130_fd_sc_hd__nor2_1 _22711_ (.A(_04834_),
    .B(_09142_),
    .Y(_02214_));
 sky130_fd_sc_hd__nor2_1 _22712_ (.A(_04843_),
    .B(_09142_),
    .Y(_02215_));
 sky130_fd_sc_hd__nor2_1 _22713_ (.A(_04852_),
    .B(_09142_),
    .Y(_02216_));
 sky130_fd_sc_hd__nor2_1 _22714_ (.A(_04860_),
    .B(_09142_),
    .Y(_02217_));
 sky130_fd_sc_hd__nand2_8 _22715_ (.A(_09825_),
    .B(_05557_),
    .Y(_09146_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_680 ();
 sky130_fd_sc_hd__nor2_1 _22717_ (.A(_05118_),
    .B(_09146_),
    .Y(_02218_));
 sky130_fd_sc_hd__nor2_1 _22718_ (.A(_05192_),
    .B(_09146_),
    .Y(_02219_));
 sky130_fd_sc_hd__nor2_1 _22719_ (.A(_05204_),
    .B(_09146_),
    .Y(_02220_));
 sky130_fd_sc_hd__nor2_1 _22720_ (.A(_05214_),
    .B(_09146_),
    .Y(_02221_));
 sky130_fd_sc_hd__nor2_1 _22721_ (.A(_05221_),
    .B(_09146_),
    .Y(_02222_));
 sky130_fd_sc_hd__nor2_1 _22722_ (.A(net1138),
    .B(_09146_),
    .Y(_02223_));
 sky130_fd_sc_hd__nor2_1 _22723_ (.A(_05238_),
    .B(_09146_),
    .Y(_02224_));
 sky130_fd_sc_hd__nor2_1 _22724_ (.A(net1140),
    .B(_09146_),
    .Y(_02225_));
 sky130_fd_sc_hd__nor2_1 _22725_ (.A(_05258_),
    .B(_09146_),
    .Y(_02226_));
 sky130_fd_sc_hd__nor2_1 _22726_ (.A(net1136),
    .B(_09146_),
    .Y(_02227_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_679 ();
 sky130_fd_sc_hd__nor2_1 _22728_ (.A(_05280_),
    .B(_09146_),
    .Y(_02228_));
 sky130_fd_sc_hd__nor2_1 _22729_ (.A(_05122_),
    .B(_09146_),
    .Y(_02229_));
 sky130_fd_sc_hd__nor2_1 _22730_ (.A(_05291_),
    .B(_09146_),
    .Y(_02230_));
 sky130_fd_sc_hd__nor2_1 _22731_ (.A(_05301_),
    .B(_09146_),
    .Y(_02231_));
 sky130_fd_sc_hd__nor2_1 _22732_ (.A(_05309_),
    .B(_09146_),
    .Y(_02232_));
 sky130_fd_sc_hd__nor2_1 _22733_ (.A(_05320_),
    .B(_09146_),
    .Y(_02233_));
 sky130_fd_sc_hd__nor2_1 _22734_ (.A(net1112),
    .B(_09146_),
    .Y(_02234_));
 sky130_fd_sc_hd__nor2_1 _22735_ (.A(_05339_),
    .B(_09146_),
    .Y(_02235_));
 sky130_fd_sc_hd__nor2_1 _22736_ (.A(net1144),
    .B(_09146_),
    .Y(_02236_));
 sky130_fd_sc_hd__nor2_1 _22737_ (.A(_05358_),
    .B(_09146_),
    .Y(_02237_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_678 ();
 sky130_fd_sc_hd__nor2_1 _22739_ (.A(net1134),
    .B(_09146_),
    .Y(_02238_));
 sky130_fd_sc_hd__nor2_1 _22740_ (.A(_05380_),
    .B(_09146_),
    .Y(_02239_));
 sky130_fd_sc_hd__nor2_1 _22741_ (.A(_05126_),
    .B(_09146_),
    .Y(_02240_));
 sky130_fd_sc_hd__nor2_1 _22742_ (.A(net1114),
    .B(_09146_),
    .Y(_02241_));
 sky130_fd_sc_hd__nor2_1 _22743_ (.A(_05430_),
    .B(_09146_),
    .Y(_02242_));
 sky130_fd_sc_hd__nor2_1 _22744_ (.A(_05132_),
    .B(_09146_),
    .Y(_02243_));
 sky130_fd_sc_hd__nor2_1 _22745_ (.A(_05140_),
    .B(_09146_),
    .Y(_02244_));
 sky130_fd_sc_hd__nor2_1 _22746_ (.A(_05149_),
    .B(_09146_),
    .Y(_02245_));
 sky130_fd_sc_hd__nor2_1 _22747_ (.A(_05157_),
    .B(_09146_),
    .Y(_02246_));
 sky130_fd_sc_hd__nor2_1 _22748_ (.A(_05166_),
    .B(_09146_),
    .Y(_02247_));
 sky130_fd_sc_hd__nor2_1 _22749_ (.A(_05173_),
    .B(_09146_),
    .Y(_02248_));
 sky130_fd_sc_hd__nor2_1 _22750_ (.A(_05183_),
    .B(_09146_),
    .Y(_02249_));
 sky130_fd_sc_hd__nand2_8 _22751_ (.A(_09771_),
    .B(_05598_),
    .Y(_09150_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_677 ();
 sky130_fd_sc_hd__nor2_1 _22753_ (.A(_04790_),
    .B(_09150_),
    .Y(_02250_));
 sky130_fd_sc_hd__nor2_1 _22754_ (.A(_04871_),
    .B(_09150_),
    .Y(_02251_));
 sky130_fd_sc_hd__nor2_1 _22755_ (.A(_04883_),
    .B(_09150_),
    .Y(_02252_));
 sky130_fd_sc_hd__nor2_1 _22756_ (.A(_04892_),
    .B(_09150_),
    .Y(_02253_));
 sky130_fd_sc_hd__nor2_1 _22757_ (.A(_04899_),
    .B(_09150_),
    .Y(_02254_));
 sky130_fd_sc_hd__nor2_1 _22758_ (.A(_04906_),
    .B(_09150_),
    .Y(_02255_));
 sky130_fd_sc_hd__nor2_1 _22759_ (.A(_04913_),
    .B(_09150_),
    .Y(_02256_));
 sky130_fd_sc_hd__nor2_1 _22760_ (.A(_04923_),
    .B(_09150_),
    .Y(_02257_));
 sky130_fd_sc_hd__nor2_1 _22761_ (.A(_04932_),
    .B(_09150_),
    .Y(_02258_));
 sky130_fd_sc_hd__nor2_1 _22762_ (.A(net1142),
    .B(_09150_),
    .Y(_02259_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_676 ();
 sky130_fd_sc_hd__nor2_1 _22764_ (.A(_04951_),
    .B(_09150_),
    .Y(_02260_));
 sky130_fd_sc_hd__nor2_1 _22765_ (.A(_04794_),
    .B(_09150_),
    .Y(_02261_));
 sky130_fd_sc_hd__nor2_1 _22766_ (.A(_04960_),
    .B(_09150_),
    .Y(_02262_));
 sky130_fd_sc_hd__nor2_1 _22767_ (.A(_04974_),
    .B(_09150_),
    .Y(_02263_));
 sky130_fd_sc_hd__nor2_1 _22768_ (.A(net1137),
    .B(_09150_),
    .Y(_02264_));
 sky130_fd_sc_hd__nor2_1 _22769_ (.A(_04990_),
    .B(_09150_),
    .Y(_02265_));
 sky130_fd_sc_hd__nor2_1 _22770_ (.A(net1128),
    .B(_09150_),
    .Y(_02266_));
 sky130_fd_sc_hd__nor2_1 _22771_ (.A(_05011_),
    .B(_09150_),
    .Y(_02267_));
 sky130_fd_sc_hd__nor2_1 _22772_ (.A(net1139),
    .B(_09150_),
    .Y(_02268_));
 sky130_fd_sc_hd__nor2_1 _22773_ (.A(_05029_),
    .B(_09150_),
    .Y(_02269_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_675 ();
 sky130_fd_sc_hd__nor2_1 _22775_ (.A(net1135),
    .B(_09150_),
    .Y(_02270_));
 sky130_fd_sc_hd__nor2_1 _22776_ (.A(_05044_),
    .B(_09150_),
    .Y(_02271_));
 sky130_fd_sc_hd__nor2_1 _22777_ (.A(_04801_),
    .B(_09150_),
    .Y(_02272_));
 sky130_fd_sc_hd__nor2_1 _22778_ (.A(_05060_),
    .B(_09150_),
    .Y(_02273_));
 sky130_fd_sc_hd__nor2_1 _22779_ (.A(_08895_),
    .B(_09150_),
    .Y(_02274_));
 sky130_fd_sc_hd__nor2_1 _22780_ (.A(_04808_),
    .B(_09150_),
    .Y(_02275_));
 sky130_fd_sc_hd__nor2_1 _22781_ (.A(_04817_),
    .B(_09150_),
    .Y(_02276_));
 sky130_fd_sc_hd__nor2_1 _22782_ (.A(_04826_),
    .B(_09150_),
    .Y(_02277_));
 sky130_fd_sc_hd__nor2_1 _22783_ (.A(_04834_),
    .B(_09150_),
    .Y(_02278_));
 sky130_fd_sc_hd__nor2_1 _22784_ (.A(_04843_),
    .B(_09150_),
    .Y(_02279_));
 sky130_fd_sc_hd__nor2_1 _22785_ (.A(_04852_),
    .B(_09150_),
    .Y(_02280_));
 sky130_fd_sc_hd__nor2_1 _22786_ (.A(_04860_),
    .B(_09150_),
    .Y(_02281_));
 sky130_fd_sc_hd__or3_4 _22787_ (.A(net1039),
    .B(_09816_),
    .C(_09793_),
    .X(_09154_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_673 ();
 sky130_fd_sc_hd__nor2_1 _22790_ (.A(_05118_),
    .B(_09154_),
    .Y(_02282_));
 sky130_fd_sc_hd__nor2_1 _22791_ (.A(_05192_),
    .B(_09154_),
    .Y(_02283_));
 sky130_fd_sc_hd__nor2_1 _22792_ (.A(_05204_),
    .B(_09154_),
    .Y(_02284_));
 sky130_fd_sc_hd__nor2_1 _22793_ (.A(_05214_),
    .B(_09154_),
    .Y(_02285_));
 sky130_fd_sc_hd__nor2_1 _22794_ (.A(_05221_),
    .B(_09154_),
    .Y(_02286_));
 sky130_fd_sc_hd__nor2_1 _22795_ (.A(_05228_),
    .B(_09154_),
    .Y(_02287_));
 sky130_fd_sc_hd__nor2_1 _22796_ (.A(_05238_),
    .B(_09154_),
    .Y(_02288_));
 sky130_fd_sc_hd__nor2_1 _22797_ (.A(net1140),
    .B(_09154_),
    .Y(_02289_));
 sky130_fd_sc_hd__nor2_1 _22798_ (.A(_05258_),
    .B(_09154_),
    .Y(_02290_));
 sky130_fd_sc_hd__nor2_1 _22799_ (.A(net1136),
    .B(_09154_),
    .Y(_02291_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_672 ();
 sky130_fd_sc_hd__nor2_1 _22801_ (.A(_05280_),
    .B(_09154_),
    .Y(_02292_));
 sky130_fd_sc_hd__nor2_1 _22802_ (.A(_05122_),
    .B(_09154_),
    .Y(_02293_));
 sky130_fd_sc_hd__nor2_1 _22803_ (.A(_05291_),
    .B(_09154_),
    .Y(_02294_));
 sky130_fd_sc_hd__nor2_1 _22804_ (.A(_05301_),
    .B(_09154_),
    .Y(_02295_));
 sky130_fd_sc_hd__nor2_1 _22805_ (.A(_05309_),
    .B(_09154_),
    .Y(_02296_));
 sky130_fd_sc_hd__nor2_1 _22806_ (.A(_05320_),
    .B(_09154_),
    .Y(_02297_));
 sky130_fd_sc_hd__nor2_1 _22807_ (.A(net1112),
    .B(_09154_),
    .Y(_02298_));
 sky130_fd_sc_hd__nor2_1 _22808_ (.A(_05339_),
    .B(_09154_),
    .Y(_02299_));
 sky130_fd_sc_hd__nor2_1 _22809_ (.A(_05347_),
    .B(_09154_),
    .Y(_02300_));
 sky130_fd_sc_hd__nor2_1 _22810_ (.A(_05358_),
    .B(_09154_),
    .Y(_02301_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_671 ();
 sky130_fd_sc_hd__nor2_1 _22812_ (.A(net1141),
    .B(_09154_),
    .Y(_02302_));
 sky130_fd_sc_hd__nor2_1 _22813_ (.A(_05380_),
    .B(_09154_),
    .Y(_02303_));
 sky130_fd_sc_hd__nor2_1 _22814_ (.A(_05126_),
    .B(_09154_),
    .Y(_02304_));
 sky130_fd_sc_hd__nor2_1 _22815_ (.A(net1143),
    .B(_09154_),
    .Y(_02305_));
 sky130_fd_sc_hd__nor2_1 _22816_ (.A(_05430_),
    .B(_09154_),
    .Y(_02306_));
 sky130_fd_sc_hd__nor2_1 _22817_ (.A(_05132_),
    .B(_09154_),
    .Y(_02307_));
 sky130_fd_sc_hd__nor2_1 _22818_ (.A(_05140_),
    .B(_09154_),
    .Y(_02308_));
 sky130_fd_sc_hd__nor2_1 _22819_ (.A(_05149_),
    .B(_09154_),
    .Y(_02309_));
 sky130_fd_sc_hd__nor2_1 _22820_ (.A(_05157_),
    .B(_09154_),
    .Y(_02310_));
 sky130_fd_sc_hd__nor2_1 _22821_ (.A(_05166_),
    .B(_09154_),
    .Y(_02311_));
 sky130_fd_sc_hd__nor2_1 _22822_ (.A(_05173_),
    .B(_09154_),
    .Y(_02312_));
 sky130_fd_sc_hd__nor2_1 _22823_ (.A(_05183_),
    .B(_09154_),
    .Y(_02313_));
 sky130_fd_sc_hd__nand2_8 _22824_ (.A(_09778_),
    .B(_04784_),
    .Y(_09159_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_670 ();
 sky130_fd_sc_hd__nor2_1 _22826_ (.A(_04790_),
    .B(_09159_),
    .Y(_02314_));
 sky130_fd_sc_hd__nor2_1 _22827_ (.A(_04871_),
    .B(_09159_),
    .Y(_02315_));
 sky130_fd_sc_hd__nor2_1 _22828_ (.A(_04883_),
    .B(_09159_),
    .Y(_02316_));
 sky130_fd_sc_hd__nor2_1 _22829_ (.A(_04892_),
    .B(_09159_),
    .Y(_02317_));
 sky130_fd_sc_hd__nor2_1 _22830_ (.A(_04899_),
    .B(_09159_),
    .Y(_02318_));
 sky130_fd_sc_hd__nor2_1 _22831_ (.A(_04906_),
    .B(_09159_),
    .Y(_02319_));
 sky130_fd_sc_hd__nor2_1 _22832_ (.A(_04913_),
    .B(_09159_),
    .Y(_02320_));
 sky130_fd_sc_hd__nor2_1 _22833_ (.A(_04923_),
    .B(_09159_),
    .Y(_02321_));
 sky130_fd_sc_hd__nor2_1 _22834_ (.A(_04932_),
    .B(_09159_),
    .Y(_02322_));
 sky130_fd_sc_hd__nor2_1 _22835_ (.A(net1142),
    .B(_09159_),
    .Y(_02323_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_669 ();
 sky130_fd_sc_hd__nor2_1 _22837_ (.A(_04951_),
    .B(_09159_),
    .Y(_02324_));
 sky130_fd_sc_hd__nor2_1 _22838_ (.A(_04794_),
    .B(_09159_),
    .Y(_02325_));
 sky130_fd_sc_hd__nor2_1 _22839_ (.A(_04960_),
    .B(_09159_),
    .Y(_02326_));
 sky130_fd_sc_hd__nor2_1 _22840_ (.A(_04974_),
    .B(_09159_),
    .Y(_02327_));
 sky130_fd_sc_hd__nor2_1 _22841_ (.A(net1137),
    .B(_09159_),
    .Y(_02328_));
 sky130_fd_sc_hd__nor2_1 _22842_ (.A(_04990_),
    .B(_09159_),
    .Y(_02329_));
 sky130_fd_sc_hd__nor2_1 _22843_ (.A(_05000_),
    .B(_09159_),
    .Y(_02330_));
 sky130_fd_sc_hd__nor2_1 _22844_ (.A(_05011_),
    .B(_09159_),
    .Y(_02331_));
 sky130_fd_sc_hd__nor2_1 _22845_ (.A(net1139),
    .B(_09159_),
    .Y(_02332_));
 sky130_fd_sc_hd__nor2_1 _22846_ (.A(_05029_),
    .B(_09159_),
    .Y(_02333_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_668 ();
 sky130_fd_sc_hd__nor2_1 _22848_ (.A(net1135),
    .B(_09159_),
    .Y(_02334_));
 sky130_fd_sc_hd__nor2_1 _22849_ (.A(_05044_),
    .B(_09159_),
    .Y(_02335_));
 sky130_fd_sc_hd__nor2_1 _22850_ (.A(_04801_),
    .B(_09159_),
    .Y(_02336_));
 sky130_fd_sc_hd__nor2_1 _22851_ (.A(_05060_),
    .B(_09159_),
    .Y(_02337_));
 sky130_fd_sc_hd__nor2_1 _22852_ (.A(_08895_),
    .B(_09159_),
    .Y(_02338_));
 sky130_fd_sc_hd__nor2_1 _22853_ (.A(_04808_),
    .B(_09159_),
    .Y(_02339_));
 sky130_fd_sc_hd__nor2_1 _22854_ (.A(_04817_),
    .B(_09159_),
    .Y(_02340_));
 sky130_fd_sc_hd__nor2_1 _22855_ (.A(_04826_),
    .B(_09159_),
    .Y(_02341_));
 sky130_fd_sc_hd__nor2_1 _22856_ (.A(_04834_),
    .B(_09159_),
    .Y(_02342_));
 sky130_fd_sc_hd__nor2_1 _22857_ (.A(_04843_),
    .B(_09159_),
    .Y(_02343_));
 sky130_fd_sc_hd__nor2_1 _22858_ (.A(_04852_),
    .B(_09159_),
    .Y(_02344_));
 sky130_fd_sc_hd__nor2_1 _22859_ (.A(_04860_),
    .B(_09159_),
    .Y(_02345_));
 sky130_fd_sc_hd__nand2_8 _22860_ (.A(_09830_),
    .B(_05115_),
    .Y(_09163_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_667 ();
 sky130_fd_sc_hd__nor2_1 _22862_ (.A(_05118_),
    .B(_09163_),
    .Y(_02346_));
 sky130_fd_sc_hd__nor2_1 _22863_ (.A(_05192_),
    .B(_09163_),
    .Y(_02347_));
 sky130_fd_sc_hd__nor2_1 _22864_ (.A(_05204_),
    .B(_09163_),
    .Y(_02348_));
 sky130_fd_sc_hd__nor2_1 _22865_ (.A(_05214_),
    .B(_09163_),
    .Y(_02349_));
 sky130_fd_sc_hd__nor2_1 _22866_ (.A(_05221_),
    .B(_09163_),
    .Y(_02350_));
 sky130_fd_sc_hd__nor2_1 _22867_ (.A(net1138),
    .B(_09163_),
    .Y(_02351_));
 sky130_fd_sc_hd__nor2_1 _22868_ (.A(_05238_),
    .B(_09163_),
    .Y(_02352_));
 sky130_fd_sc_hd__nor2_1 _22869_ (.A(net1140),
    .B(_09163_),
    .Y(_02353_));
 sky130_fd_sc_hd__nor2_1 _22870_ (.A(_05258_),
    .B(_09163_),
    .Y(_02354_));
 sky130_fd_sc_hd__nor2_1 _22871_ (.A(_05267_),
    .B(_09163_),
    .Y(_02355_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_666 ();
 sky130_fd_sc_hd__nor2_1 _22873_ (.A(_05280_),
    .B(_09163_),
    .Y(_02356_));
 sky130_fd_sc_hd__nor2_1 _22874_ (.A(_05122_),
    .B(_09163_),
    .Y(_02357_));
 sky130_fd_sc_hd__nor2_1 _22875_ (.A(_05291_),
    .B(_09163_),
    .Y(_02358_));
 sky130_fd_sc_hd__nor2_1 _22876_ (.A(_05301_),
    .B(_09163_),
    .Y(_02359_));
 sky130_fd_sc_hd__nor2_1 _22877_ (.A(_05309_),
    .B(_09163_),
    .Y(_02360_));
 sky130_fd_sc_hd__nor2_1 _22878_ (.A(_05320_),
    .B(_09163_),
    .Y(_02361_));
 sky130_fd_sc_hd__nor2_1 _22879_ (.A(net1112),
    .B(_09163_),
    .Y(_02362_));
 sky130_fd_sc_hd__nor2_1 _22880_ (.A(_05339_),
    .B(_09163_),
    .Y(_02363_));
 sky130_fd_sc_hd__nor2_1 _22881_ (.A(_05347_),
    .B(_09163_),
    .Y(_02364_));
 sky130_fd_sc_hd__nor2_1 _22882_ (.A(_05358_),
    .B(_09163_),
    .Y(_02365_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_665 ();
 sky130_fd_sc_hd__nor2_1 _22884_ (.A(net1134),
    .B(_09163_),
    .Y(_02366_));
 sky130_fd_sc_hd__nor2_1 _22885_ (.A(_05380_),
    .B(_09163_),
    .Y(_02367_));
 sky130_fd_sc_hd__nor2_1 _22886_ (.A(_05126_),
    .B(_09163_),
    .Y(_02368_));
 sky130_fd_sc_hd__nor2_1 _22887_ (.A(net1114),
    .B(_09163_),
    .Y(_02369_));
 sky130_fd_sc_hd__nor2_1 _22888_ (.A(_05430_),
    .B(_09163_),
    .Y(_02370_));
 sky130_fd_sc_hd__nor2_1 _22889_ (.A(_05132_),
    .B(_09163_),
    .Y(_02371_));
 sky130_fd_sc_hd__nor2_1 _22890_ (.A(_05140_),
    .B(_09163_),
    .Y(_02372_));
 sky130_fd_sc_hd__nor2_1 _22891_ (.A(_05149_),
    .B(_09163_),
    .Y(_02373_));
 sky130_fd_sc_hd__nor2_1 _22892_ (.A(_05157_),
    .B(_09163_),
    .Y(_02374_));
 sky130_fd_sc_hd__nor2_1 _22893_ (.A(_05166_),
    .B(_09163_),
    .Y(_02375_));
 sky130_fd_sc_hd__nor2_1 _22894_ (.A(_05173_),
    .B(_09163_),
    .Y(_02376_));
 sky130_fd_sc_hd__nor2_1 _22895_ (.A(_05183_),
    .B(_09163_),
    .Y(_02377_));
 sky130_fd_sc_hd__nand2_8 _22896_ (.A(_09778_),
    .B(_05433_),
    .Y(_09167_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_664 ();
 sky130_fd_sc_hd__nor2_1 _22898_ (.A(_04790_),
    .B(_09167_),
    .Y(_02378_));
 sky130_fd_sc_hd__nor2_1 _22899_ (.A(_04871_),
    .B(_09167_),
    .Y(_02379_));
 sky130_fd_sc_hd__nor2_1 _22900_ (.A(_04883_),
    .B(_09167_),
    .Y(_02380_));
 sky130_fd_sc_hd__nor2_1 _22901_ (.A(_04892_),
    .B(_09167_),
    .Y(_02381_));
 sky130_fd_sc_hd__nor2_1 _22902_ (.A(_04899_),
    .B(_09167_),
    .Y(_02382_));
 sky130_fd_sc_hd__nor2_1 _22903_ (.A(_04906_),
    .B(_09167_),
    .Y(_02383_));
 sky130_fd_sc_hd__nor2_1 _22904_ (.A(_04913_),
    .B(_09167_),
    .Y(_02384_));
 sky130_fd_sc_hd__nor2_1 _22905_ (.A(_04923_),
    .B(_09167_),
    .Y(_02385_));
 sky130_fd_sc_hd__nor2_1 _22906_ (.A(_04932_),
    .B(_09167_),
    .Y(_02386_));
 sky130_fd_sc_hd__nor2_1 _22907_ (.A(net1142),
    .B(_09167_),
    .Y(_02387_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_663 ();
 sky130_fd_sc_hd__nor2_1 _22909_ (.A(_04951_),
    .B(_09167_),
    .Y(_02388_));
 sky130_fd_sc_hd__nor2_1 _22910_ (.A(_04794_),
    .B(_09167_),
    .Y(_02389_));
 sky130_fd_sc_hd__nor2_1 _22911_ (.A(_04960_),
    .B(_09167_),
    .Y(_02390_));
 sky130_fd_sc_hd__nor2_1 _22912_ (.A(_04974_),
    .B(_09167_),
    .Y(_02391_));
 sky130_fd_sc_hd__nor2_1 _22913_ (.A(net1137),
    .B(_09167_),
    .Y(_02392_));
 sky130_fd_sc_hd__nor2_1 _22914_ (.A(_04990_),
    .B(_09167_),
    .Y(_02393_));
 sky130_fd_sc_hd__nor2_1 _22915_ (.A(net1128),
    .B(_09167_),
    .Y(_02394_));
 sky130_fd_sc_hd__nor2_1 _22916_ (.A(_05011_),
    .B(_09167_),
    .Y(_02395_));
 sky130_fd_sc_hd__nor2_1 _22917_ (.A(_05020_),
    .B(_09167_),
    .Y(_02396_));
 sky130_fd_sc_hd__nor2_1 _22918_ (.A(_05029_),
    .B(_09167_),
    .Y(_02397_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_662 ();
 sky130_fd_sc_hd__nor2_1 _22920_ (.A(net1135),
    .B(_09167_),
    .Y(_02398_));
 sky130_fd_sc_hd__nor2_1 _22921_ (.A(_05044_),
    .B(_09167_),
    .Y(_02399_));
 sky130_fd_sc_hd__nor2_1 _22922_ (.A(_04801_),
    .B(_09167_),
    .Y(_02400_));
 sky130_fd_sc_hd__nor2_1 _22923_ (.A(_05060_),
    .B(_09167_),
    .Y(_02401_));
 sky130_fd_sc_hd__nor2_1 _22924_ (.A(_08895_),
    .B(_09167_),
    .Y(_02402_));
 sky130_fd_sc_hd__nor2_1 _22925_ (.A(_04808_),
    .B(_09167_),
    .Y(_02403_));
 sky130_fd_sc_hd__nor2_1 _22926_ (.A(_04817_),
    .B(_09167_),
    .Y(_02404_));
 sky130_fd_sc_hd__nor2_1 _22927_ (.A(_04826_),
    .B(_09167_),
    .Y(_02405_));
 sky130_fd_sc_hd__nor2_1 _22928_ (.A(_04834_),
    .B(_09167_),
    .Y(_02406_));
 sky130_fd_sc_hd__nor2_1 _22929_ (.A(_04843_),
    .B(_09167_),
    .Y(_02407_));
 sky130_fd_sc_hd__nor2_1 _22930_ (.A(_04852_),
    .B(_09167_),
    .Y(_02408_));
 sky130_fd_sc_hd__nor2_1 _22931_ (.A(_04860_),
    .B(_09167_),
    .Y(_02409_));
 sky130_fd_sc_hd__nand2_8 _22932_ (.A(_09830_),
    .B(_05474_),
    .Y(_09171_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_661 ();
 sky130_fd_sc_hd__nor2_1 _22934_ (.A(_05118_),
    .B(_09171_),
    .Y(_02410_));
 sky130_fd_sc_hd__nor2_1 _22935_ (.A(_05192_),
    .B(_09171_),
    .Y(_02411_));
 sky130_fd_sc_hd__nor2_1 _22936_ (.A(_05204_),
    .B(_09171_),
    .Y(_02412_));
 sky130_fd_sc_hd__nor2_1 _22937_ (.A(_05214_),
    .B(_09171_),
    .Y(_02413_));
 sky130_fd_sc_hd__nor2_1 _22938_ (.A(_05221_),
    .B(_09171_),
    .Y(_02414_));
 sky130_fd_sc_hd__nor2_1 _22939_ (.A(_05228_),
    .B(_09171_),
    .Y(_02415_));
 sky130_fd_sc_hd__nor2_1 _22940_ (.A(_05238_),
    .B(_09171_),
    .Y(_02416_));
 sky130_fd_sc_hd__nor2_1 _22941_ (.A(net1140),
    .B(_09171_),
    .Y(_02417_));
 sky130_fd_sc_hd__nor2_1 _22942_ (.A(_05258_),
    .B(_09171_),
    .Y(_02418_));
 sky130_fd_sc_hd__nor2_1 _22943_ (.A(net1136),
    .B(_09171_),
    .Y(_02419_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_660 ();
 sky130_fd_sc_hd__nor2_1 _22945_ (.A(_05280_),
    .B(_09171_),
    .Y(_02420_));
 sky130_fd_sc_hd__nor2_1 _22946_ (.A(_05122_),
    .B(_09171_),
    .Y(_02421_));
 sky130_fd_sc_hd__nor2_1 _22947_ (.A(_05291_),
    .B(_09171_),
    .Y(_02422_));
 sky130_fd_sc_hd__nor2_1 _22948_ (.A(_05301_),
    .B(_09171_),
    .Y(_02423_));
 sky130_fd_sc_hd__nor2_1 _22949_ (.A(_05309_),
    .B(_09171_),
    .Y(_02424_));
 sky130_fd_sc_hd__nor2_1 _22950_ (.A(_05320_),
    .B(_09171_),
    .Y(_02425_));
 sky130_fd_sc_hd__nor2_1 _22951_ (.A(net1112),
    .B(_09171_),
    .Y(_02426_));
 sky130_fd_sc_hd__nor2_1 _22952_ (.A(_05339_),
    .B(_09171_),
    .Y(_02427_));
 sky130_fd_sc_hd__nor2_1 _22953_ (.A(_05347_),
    .B(_09171_),
    .Y(_02428_));
 sky130_fd_sc_hd__nor2_1 _22954_ (.A(_05358_),
    .B(_09171_),
    .Y(_02429_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_659 ();
 sky130_fd_sc_hd__nor2_1 _22956_ (.A(net1134),
    .B(_09171_),
    .Y(_02430_));
 sky130_fd_sc_hd__nor2_1 _22957_ (.A(_05380_),
    .B(_09171_),
    .Y(_02431_));
 sky130_fd_sc_hd__nor2_1 _22958_ (.A(_05126_),
    .B(_09171_),
    .Y(_02432_));
 sky130_fd_sc_hd__nor2_1 _22959_ (.A(net1143),
    .B(_09171_),
    .Y(_02433_));
 sky130_fd_sc_hd__nor2_1 _22960_ (.A(_05430_),
    .B(_09171_),
    .Y(_02434_));
 sky130_fd_sc_hd__nor2_1 _22961_ (.A(_05132_),
    .B(_09171_),
    .Y(_02435_));
 sky130_fd_sc_hd__nor2_1 _22962_ (.A(_05140_),
    .B(_09171_),
    .Y(_02436_));
 sky130_fd_sc_hd__nor2_1 _22963_ (.A(_05149_),
    .B(_09171_),
    .Y(_02437_));
 sky130_fd_sc_hd__nor2_1 _22964_ (.A(_05157_),
    .B(_09171_),
    .Y(_02438_));
 sky130_fd_sc_hd__nor2_1 _22965_ (.A(_05166_),
    .B(_09171_),
    .Y(_02439_));
 sky130_fd_sc_hd__nor2_1 _22966_ (.A(_05173_),
    .B(_09171_),
    .Y(_02440_));
 sky130_fd_sc_hd__nor2_1 _22967_ (.A(_05183_),
    .B(_09171_),
    .Y(_02441_));
 sky130_fd_sc_hd__nand2_8 _22968_ (.A(_09778_),
    .B(_05516_),
    .Y(_09175_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_658 ();
 sky130_fd_sc_hd__nor2_1 _22970_ (.A(_04790_),
    .B(_09175_),
    .Y(_02442_));
 sky130_fd_sc_hd__nor2_1 _22971_ (.A(_04871_),
    .B(_09175_),
    .Y(_02443_));
 sky130_fd_sc_hd__nor2_1 _22972_ (.A(_04883_),
    .B(_09175_),
    .Y(_02444_));
 sky130_fd_sc_hd__nor2_1 _22973_ (.A(_04892_),
    .B(_09175_),
    .Y(_02445_));
 sky130_fd_sc_hd__nor2_1 _22974_ (.A(_04899_),
    .B(_09175_),
    .Y(_02446_));
 sky130_fd_sc_hd__nor2_1 _22975_ (.A(_04906_),
    .B(_09175_),
    .Y(_02447_));
 sky130_fd_sc_hd__nor2_1 _22976_ (.A(_04913_),
    .B(_09175_),
    .Y(_02448_));
 sky130_fd_sc_hd__nor2_1 _22977_ (.A(_04923_),
    .B(_09175_),
    .Y(_02449_));
 sky130_fd_sc_hd__nor2_1 _22978_ (.A(_04932_),
    .B(_09175_),
    .Y(_02450_));
 sky130_fd_sc_hd__nor2_1 _22979_ (.A(_04939_),
    .B(_09175_),
    .Y(_02451_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_657 ();
 sky130_fd_sc_hd__nor2_1 _22981_ (.A(_04951_),
    .B(_09175_),
    .Y(_02452_));
 sky130_fd_sc_hd__nor2_1 _22982_ (.A(_04794_),
    .B(_09175_),
    .Y(_02453_));
 sky130_fd_sc_hd__nor2_1 _22983_ (.A(_04960_),
    .B(_09175_),
    .Y(_02454_));
 sky130_fd_sc_hd__nor2_1 _22984_ (.A(_04974_),
    .B(_09175_),
    .Y(_02455_));
 sky130_fd_sc_hd__nor2_1 _22985_ (.A(net1137),
    .B(_09175_),
    .Y(_02456_));
 sky130_fd_sc_hd__nor2_1 _22986_ (.A(_04990_),
    .B(_09175_),
    .Y(_02457_));
 sky130_fd_sc_hd__nor2_1 _22987_ (.A(net1128),
    .B(_09175_),
    .Y(_02458_));
 sky130_fd_sc_hd__nor2_1 _22988_ (.A(_05011_),
    .B(_09175_),
    .Y(_02459_));
 sky130_fd_sc_hd__nor2_1 _22989_ (.A(net1139),
    .B(_09175_),
    .Y(_02460_));
 sky130_fd_sc_hd__nor2_1 _22990_ (.A(_05029_),
    .B(_09175_),
    .Y(_02461_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_656 ();
 sky130_fd_sc_hd__nor2_1 _22992_ (.A(net1135),
    .B(_09175_),
    .Y(_02462_));
 sky130_fd_sc_hd__nor2_1 _22993_ (.A(_05044_),
    .B(_09175_),
    .Y(_02463_));
 sky130_fd_sc_hd__nor2_1 _22994_ (.A(_04801_),
    .B(_09175_),
    .Y(_02464_));
 sky130_fd_sc_hd__nor2_1 _22995_ (.A(_05060_),
    .B(_09175_),
    .Y(_02465_));
 sky130_fd_sc_hd__nor2_1 _22996_ (.A(_08895_),
    .B(_09175_),
    .Y(_02466_));
 sky130_fd_sc_hd__nor2_1 _22997_ (.A(_04808_),
    .B(_09175_),
    .Y(_02467_));
 sky130_fd_sc_hd__nor2_1 _22998_ (.A(_04817_),
    .B(_09175_),
    .Y(_02468_));
 sky130_fd_sc_hd__nor2_1 _22999_ (.A(_04826_),
    .B(_09175_),
    .Y(_02469_));
 sky130_fd_sc_hd__nor2_1 _23000_ (.A(_04834_),
    .B(_09175_),
    .Y(_02470_));
 sky130_fd_sc_hd__nor2_1 _23001_ (.A(_04843_),
    .B(_09175_),
    .Y(_02471_));
 sky130_fd_sc_hd__nor2_1 _23002_ (.A(_04852_),
    .B(_09175_),
    .Y(_02472_));
 sky130_fd_sc_hd__nor2_1 _23003_ (.A(_04860_),
    .B(_09175_),
    .Y(_02473_));
 sky130_fd_sc_hd__nand2_8 _23004_ (.A(_09830_),
    .B(_05557_),
    .Y(_09179_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_655 ();
 sky130_fd_sc_hd__nor2_1 _23006_ (.A(_05118_),
    .B(_09179_),
    .Y(_02474_));
 sky130_fd_sc_hd__nor2_1 _23007_ (.A(_05192_),
    .B(_09179_),
    .Y(_02475_));
 sky130_fd_sc_hd__nor2_1 _23008_ (.A(_05204_),
    .B(_09179_),
    .Y(_02476_));
 sky130_fd_sc_hd__nor2_1 _23009_ (.A(_05214_),
    .B(_09179_),
    .Y(_02477_));
 sky130_fd_sc_hd__nor2_1 _23010_ (.A(_05221_),
    .B(_09179_),
    .Y(_02478_));
 sky130_fd_sc_hd__nor2_1 _23011_ (.A(net1138),
    .B(_09179_),
    .Y(_02479_));
 sky130_fd_sc_hd__nor2_1 _23012_ (.A(_05238_),
    .B(_09179_),
    .Y(_02480_));
 sky130_fd_sc_hd__nor2_1 _23013_ (.A(net1140),
    .B(_09179_),
    .Y(_02481_));
 sky130_fd_sc_hd__nor2_1 _23014_ (.A(_05258_),
    .B(_09179_),
    .Y(_02482_));
 sky130_fd_sc_hd__nor2_1 _23015_ (.A(net1136),
    .B(_09179_),
    .Y(_02483_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_654 ();
 sky130_fd_sc_hd__nor2_1 _23017_ (.A(_05280_),
    .B(_09179_),
    .Y(_02484_));
 sky130_fd_sc_hd__nor2_1 _23018_ (.A(_05122_),
    .B(_09179_),
    .Y(_02485_));
 sky130_fd_sc_hd__nor2_1 _23019_ (.A(_05291_),
    .B(_09179_),
    .Y(_02486_));
 sky130_fd_sc_hd__nor2_1 _23020_ (.A(_05301_),
    .B(_09179_),
    .Y(_02487_));
 sky130_fd_sc_hd__nor2_1 _23021_ (.A(_05309_),
    .B(_09179_),
    .Y(_02488_));
 sky130_fd_sc_hd__nor2_1 _23022_ (.A(_05320_),
    .B(_09179_),
    .Y(_02489_));
 sky130_fd_sc_hd__nor2_1 _23023_ (.A(net1112),
    .B(_09179_),
    .Y(_02490_));
 sky130_fd_sc_hd__nor2_1 _23024_ (.A(_05339_),
    .B(_09179_),
    .Y(_02491_));
 sky130_fd_sc_hd__nor2_1 _23025_ (.A(net1144),
    .B(_09179_),
    .Y(_02492_));
 sky130_fd_sc_hd__nor2_1 _23026_ (.A(_05358_),
    .B(_09179_),
    .Y(_02493_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_653 ();
 sky130_fd_sc_hd__nor2_1 _23028_ (.A(net1134),
    .B(_09179_),
    .Y(_02494_));
 sky130_fd_sc_hd__nor2_1 _23029_ (.A(_05380_),
    .B(_09179_),
    .Y(_02495_));
 sky130_fd_sc_hd__nor2_1 _23030_ (.A(_05126_),
    .B(_09179_),
    .Y(_02496_));
 sky130_fd_sc_hd__nor2_1 _23031_ (.A(net1143),
    .B(_09179_),
    .Y(_02497_));
 sky130_fd_sc_hd__nor2_1 _23032_ (.A(_05430_),
    .B(_09179_),
    .Y(_02498_));
 sky130_fd_sc_hd__nor2_1 _23033_ (.A(_05132_),
    .B(_09179_),
    .Y(_02499_));
 sky130_fd_sc_hd__nor2_1 _23034_ (.A(_05140_),
    .B(_09179_),
    .Y(_02500_));
 sky130_fd_sc_hd__nor2_1 _23035_ (.A(_05149_),
    .B(_09179_),
    .Y(_02501_));
 sky130_fd_sc_hd__nor2_1 _23036_ (.A(_05157_),
    .B(_09179_),
    .Y(_02502_));
 sky130_fd_sc_hd__nor2_1 _23037_ (.A(_05166_),
    .B(_09179_),
    .Y(_02503_));
 sky130_fd_sc_hd__nor2_1 _23038_ (.A(_05173_),
    .B(_09179_),
    .Y(_02504_));
 sky130_fd_sc_hd__nor2_1 _23039_ (.A(_05183_),
    .B(_09179_),
    .Y(_02505_));
 sky130_fd_sc_hd__nand2_8 _23040_ (.A(_09778_),
    .B(_05598_),
    .Y(_09183_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_652 ();
 sky130_fd_sc_hd__nor2_1 _23042_ (.A(_04790_),
    .B(_09183_),
    .Y(_02506_));
 sky130_fd_sc_hd__nor2_1 _23043_ (.A(_04871_),
    .B(_09183_),
    .Y(_02507_));
 sky130_fd_sc_hd__nor2_1 _23044_ (.A(_04883_),
    .B(_09183_),
    .Y(_02508_));
 sky130_fd_sc_hd__nor2_1 _23045_ (.A(_04892_),
    .B(_09183_),
    .Y(_02509_));
 sky130_fd_sc_hd__nor2_1 _23046_ (.A(_04899_),
    .B(_09183_),
    .Y(_02510_));
 sky130_fd_sc_hd__nor2_1 _23047_ (.A(_04906_),
    .B(_09183_),
    .Y(_02511_));
 sky130_fd_sc_hd__nor2_1 _23048_ (.A(_04913_),
    .B(_09183_),
    .Y(_02512_));
 sky130_fd_sc_hd__nor2_1 _23049_ (.A(_04923_),
    .B(_09183_),
    .Y(_02513_));
 sky130_fd_sc_hd__nor2_1 _23050_ (.A(_04932_),
    .B(_09183_),
    .Y(_02514_));
 sky130_fd_sc_hd__nor2_1 _23051_ (.A(net1142),
    .B(_09183_),
    .Y(_02515_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_651 ();
 sky130_fd_sc_hd__nor2_1 _23053_ (.A(_04951_),
    .B(_09183_),
    .Y(_02516_));
 sky130_fd_sc_hd__nor2_1 _23054_ (.A(_04794_),
    .B(_09183_),
    .Y(_02517_));
 sky130_fd_sc_hd__nor2_1 _23055_ (.A(_04960_),
    .B(_09183_),
    .Y(_02518_));
 sky130_fd_sc_hd__nor2_1 _23056_ (.A(_04974_),
    .B(_09183_),
    .Y(_02519_));
 sky130_fd_sc_hd__nor2_1 _23057_ (.A(net1137),
    .B(_09183_),
    .Y(_02520_));
 sky130_fd_sc_hd__nor2_1 _23058_ (.A(_04990_),
    .B(_09183_),
    .Y(_02521_));
 sky130_fd_sc_hd__nor2_1 _23059_ (.A(net1128),
    .B(_09183_),
    .Y(_02522_));
 sky130_fd_sc_hd__nor2_1 _23060_ (.A(_05011_),
    .B(_09183_),
    .Y(_02523_));
 sky130_fd_sc_hd__nor2_1 _23061_ (.A(_05020_),
    .B(_09183_),
    .Y(_02524_));
 sky130_fd_sc_hd__nor2_1 _23062_ (.A(_05029_),
    .B(_09183_),
    .Y(_02525_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_650 ();
 sky130_fd_sc_hd__nor2_1 _23064_ (.A(_05035_),
    .B(_09183_),
    .Y(_02526_));
 sky130_fd_sc_hd__nor2_1 _23065_ (.A(_05044_),
    .B(_09183_),
    .Y(_02527_));
 sky130_fd_sc_hd__nor2_1 _23066_ (.A(_04801_),
    .B(_09183_),
    .Y(_02528_));
 sky130_fd_sc_hd__nor2_1 _23067_ (.A(_05060_),
    .B(_09183_),
    .Y(_02529_));
 sky130_fd_sc_hd__nor2_1 _23068_ (.A(_08895_),
    .B(_09183_),
    .Y(_02530_));
 sky130_fd_sc_hd__nor2_1 _23069_ (.A(_04808_),
    .B(_09183_),
    .Y(_02531_));
 sky130_fd_sc_hd__nor2_1 _23070_ (.A(_04817_),
    .B(_09183_),
    .Y(_02532_));
 sky130_fd_sc_hd__nor2_1 _23071_ (.A(_04826_),
    .B(_09183_),
    .Y(_02533_));
 sky130_fd_sc_hd__nor2_1 _23072_ (.A(_04834_),
    .B(_09183_),
    .Y(_02534_));
 sky130_fd_sc_hd__nor2_1 _23073_ (.A(_04843_),
    .B(_09183_),
    .Y(_02535_));
 sky130_fd_sc_hd__nor2_1 _23074_ (.A(_04852_),
    .B(_09183_),
    .Y(_02536_));
 sky130_fd_sc_hd__nor2_1 _23075_ (.A(_04860_),
    .B(_09183_),
    .Y(_02537_));
 sky130_fd_sc_hd__nand2b_4 _23076_ (.A_N(_09726_),
    .B(_09731_),
    .Y(_09187_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_649 ();
 sky130_fd_sc_hd__nor2_1 _23078_ (.A(_05118_),
    .B(_09187_),
    .Y(_02538_));
 sky130_fd_sc_hd__nor2_1 _23079_ (.A(_05192_),
    .B(_09187_),
    .Y(_02539_));
 sky130_fd_sc_hd__nor2_1 _23080_ (.A(_05204_),
    .B(_09187_),
    .Y(_02540_));
 sky130_fd_sc_hd__nor2_1 _23081_ (.A(_05214_),
    .B(_09187_),
    .Y(_02541_));
 sky130_fd_sc_hd__nor2_1 _23082_ (.A(_05221_),
    .B(_09187_),
    .Y(_02542_));
 sky130_fd_sc_hd__nor2_1 _23083_ (.A(net1138),
    .B(_09187_),
    .Y(_02543_));
 sky130_fd_sc_hd__nor2_1 _23084_ (.A(_05238_),
    .B(_09187_),
    .Y(_02544_));
 sky130_fd_sc_hd__nor2_1 _23085_ (.A(_05247_),
    .B(_09187_),
    .Y(_02545_));
 sky130_fd_sc_hd__nor2_1 _23086_ (.A(_05258_),
    .B(_09187_),
    .Y(_02546_));
 sky130_fd_sc_hd__nor2_1 _23087_ (.A(net1136),
    .B(_09187_),
    .Y(_02547_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_648 ();
 sky130_fd_sc_hd__nor2_1 _23089_ (.A(_05280_),
    .B(_09187_),
    .Y(_02548_));
 sky130_fd_sc_hd__nor2_1 _23090_ (.A(_05122_),
    .B(_09187_),
    .Y(_02549_));
 sky130_fd_sc_hd__nor2_1 _23091_ (.A(_05291_),
    .B(_09187_),
    .Y(_02550_));
 sky130_fd_sc_hd__nor2_1 _23092_ (.A(_05301_),
    .B(_09187_),
    .Y(_02551_));
 sky130_fd_sc_hd__nor2_1 _23093_ (.A(_05309_),
    .B(_09187_),
    .Y(_02552_));
 sky130_fd_sc_hd__nor2_1 _23094_ (.A(_05320_),
    .B(_09187_),
    .Y(_02553_));
 sky130_fd_sc_hd__nor2_1 _23095_ (.A(net1112),
    .B(_09187_),
    .Y(_02554_));
 sky130_fd_sc_hd__nor2_1 _23096_ (.A(_05339_),
    .B(_09187_),
    .Y(_02555_));
 sky130_fd_sc_hd__nor2_1 _23097_ (.A(net1144),
    .B(_09187_),
    .Y(_02556_));
 sky130_fd_sc_hd__nor2_1 _23098_ (.A(_05358_),
    .B(_09187_),
    .Y(_02557_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_647 ();
 sky130_fd_sc_hd__nor2_1 _23100_ (.A(net1113),
    .B(_09187_),
    .Y(_02558_));
 sky130_fd_sc_hd__nor2_1 _23101_ (.A(_05380_),
    .B(_09187_),
    .Y(_02559_));
 sky130_fd_sc_hd__nor2_1 _23102_ (.A(_05126_),
    .B(_09187_),
    .Y(_02560_));
 sky130_fd_sc_hd__nor2_1 _23103_ (.A(net1114),
    .B(_09187_),
    .Y(_02561_));
 sky130_fd_sc_hd__nor2_1 _23104_ (.A(_05430_),
    .B(_09187_),
    .Y(_02562_));
 sky130_fd_sc_hd__nor2_1 _23105_ (.A(_05132_),
    .B(_09187_),
    .Y(_02563_));
 sky130_fd_sc_hd__nor2_1 _23106_ (.A(_05140_),
    .B(_09187_),
    .Y(_02564_));
 sky130_fd_sc_hd__nor2_1 _23107_ (.A(_05149_),
    .B(_09187_),
    .Y(_02565_));
 sky130_fd_sc_hd__nor2_1 _23108_ (.A(_05157_),
    .B(_09187_),
    .Y(_02566_));
 sky130_fd_sc_hd__nor2_1 _23109_ (.A(_05166_),
    .B(_09187_),
    .Y(_02567_));
 sky130_fd_sc_hd__nor2_1 _23110_ (.A(_05173_),
    .B(_09187_),
    .Y(_02568_));
 sky130_fd_sc_hd__nor2_1 _23111_ (.A(_05183_),
    .B(_09187_),
    .Y(_02569_));
 sky130_fd_sc_hd__nor2b_4 _23112_ (.A(net340),
    .B_N(\hash.CA2.b_dash[0] ),
    .Y(\hash.CA1.d[0] ));
 sky130_fd_sc_hd__clkinv_1 _23113_ (.A(_13581_),
    .Y(_09191_));
 sky130_fd_sc_hd__clkinv_2 _23114_ (.A(_13573_),
    .Y(_09192_));
 sky130_fd_sc_hd__inv_2 _23115_ (.A(_13565_),
    .Y(_09193_));
 sky130_fd_sc_hd__inv_1 _23116_ (.A(_13557_),
    .Y(_09194_));
 sky130_fd_sc_hd__nor2b_1 _23117_ (.A(_12882_),
    .B_N(_13554_),
    .Y(_09195_));
 sky130_fd_sc_hd__o21ai_2 _23118_ (.A1(_13553_),
    .A2(_09195_),
    .B1(_13558_),
    .Y(_09196_));
 sky130_fd_sc_hd__a21boi_2 _23119_ (.A1(_09194_),
    .A2(_09196_),
    .B1_N(_13562_),
    .Y(_09197_));
 sky130_fd_sc_hd__o21ai_2 _23120_ (.A1(_13561_),
    .A2(_09197_),
    .B1(_13566_),
    .Y(_09198_));
 sky130_fd_sc_hd__a21boi_2 _23121_ (.A1(_09193_),
    .A2(_09198_),
    .B1_N(_13570_),
    .Y(_09199_));
 sky130_fd_sc_hd__o21ai_2 _23122_ (.A1(_13569_),
    .A2(_09199_),
    .B1(_13574_),
    .Y(_09200_));
 sky130_fd_sc_hd__a21boi_4 _23123_ (.A1(_09192_),
    .A2(_09200_),
    .B1_N(_13578_),
    .Y(_09201_));
 sky130_fd_sc_hd__o21ai_2 _23124_ (.A1(_13577_),
    .A2(_09201_),
    .B1(_13582_),
    .Y(_09202_));
 sky130_fd_sc_hd__a21boi_4 _23125_ (.A1(_09191_),
    .A2(_09202_),
    .B1_N(_13586_),
    .Y(_09203_));
 sky130_fd_sc_hd__nand2_1 _23126_ (.A(_09191_),
    .B(_09202_),
    .Y(_09204_));
 sky130_fd_sc_hd__nor2_1 _23127_ (.A(_13586_),
    .B(_09204_),
    .Y(_09205_));
 sky130_fd_sc_hd__nor2_2 _23128_ (.A(_09203_),
    .B(_09205_),
    .Y(\hash.CA1.p1[10] ));
 sky130_fd_sc_hd__o21a_1 _23129_ (.A1(_13582_),
    .A2(_13581_),
    .B1(_13586_),
    .X(_09206_));
 sky130_fd_sc_hd__nor2_1 _23130_ (.A(_13585_),
    .B(_09206_),
    .Y(_09207_));
 sky130_fd_sc_hd__inv_2 _23131_ (.A(_13558_),
    .Y(_09208_));
 sky130_fd_sc_hd__a21o_1 _23132_ (.A1(_14204_),
    .A2(_13550_),
    .B1(_13549_),
    .X(_09209_));
 sky130_fd_sc_hd__a21oi_2 _23133_ (.A1(_13554_),
    .A2(_09209_),
    .B1(_13553_),
    .Y(_09210_));
 sky130_fd_sc_hd__nor3_2 _23134_ (.A(_13565_),
    .B(_13561_),
    .C(_13557_),
    .Y(_09211_));
 sky130_fd_sc_hd__o21ai_2 _23135_ (.A1(_09208_),
    .A2(_09210_),
    .B1(_09211_),
    .Y(_09212_));
 sky130_fd_sc_hd__o21ai_0 _23136_ (.A1(_13562_),
    .A2(_13561_),
    .B1(_13566_),
    .Y(_09213_));
 sky130_fd_sc_hd__nand2_1 _23137_ (.A(_09193_),
    .B(_09213_),
    .Y(_09214_));
 sky130_fd_sc_hd__and3_1 _23138_ (.A(_13570_),
    .B(_13574_),
    .C(_13578_),
    .X(_09215_));
 sky130_fd_sc_hd__and3_4 _23139_ (.A(_09215_),
    .B(_09214_),
    .C(_09212_),
    .X(_09216_));
 sky130_fd_sc_hd__nand2_1 _23140_ (.A(_13574_),
    .B(_13569_),
    .Y(_09217_));
 sky130_fd_sc_hd__nand2_1 _23141_ (.A(_09192_),
    .B(_09217_),
    .Y(_09218_));
 sky130_fd_sc_hd__a21oi_1 _23142_ (.A1(_13578_),
    .A2(_09218_),
    .B1(_13577_),
    .Y(_09219_));
 sky130_fd_sc_hd__nor4b_4 _23143_ (.A(_13581_),
    .B(_13585_),
    .C(_09216_),
    .D_N(_09219_),
    .Y(_09220_));
 sky130_fd_sc_hd__nor2_2 _23144_ (.A(_09207_),
    .B(_09220_),
    .Y(_09221_));
 sky130_fd_sc_hd__xor2_1 _23145_ (.A(_13590_),
    .B(_09221_),
    .X(\hash.CA1.p1[11] ));
 sky130_fd_sc_hd__o21a_1 _23146_ (.A1(_13585_),
    .A2(_09203_),
    .B1(_13590_),
    .X(_09222_));
 sky130_fd_sc_hd__nor2_1 _23147_ (.A(_13589_),
    .B(_09222_),
    .Y(_09223_));
 sky130_fd_sc_hd__xnor2_1 _23148_ (.A(_13594_),
    .B(_09223_),
    .Y(\hash.CA1.p1[12] ));
 sky130_fd_sc_hd__a21o_4 _23149_ (.A1(_13594_),
    .A2(_13589_),
    .B1(_13593_),
    .X(_09224_));
 sky130_fd_sc_hd__and3_1 _23150_ (.A(_13590_),
    .B(_13594_),
    .C(_09221_),
    .X(_09225_));
 sky130_fd_sc_hd__nor2_1 _23151_ (.A(_09224_),
    .B(_09225_),
    .Y(_09226_));
 sky130_fd_sc_hd__xnor2_1 _23152_ (.A(_13598_),
    .B(_09226_),
    .Y(\hash.CA1.p1[13] ));
 sky130_fd_sc_hd__or3_4 _23153_ (.A(_13585_),
    .B(_13597_),
    .C(_09224_),
    .X(_09227_));
 sky130_fd_sc_hd__a211oi_1 _23154_ (.A1(_13590_),
    .A2(_13594_),
    .B1(_13597_),
    .C1(_09224_),
    .Y(_09228_));
 sky130_fd_sc_hd__nor2_1 _23155_ (.A(_13598_),
    .B(_13597_),
    .Y(_09229_));
 sky130_fd_sc_hd__nor2_1 _23156_ (.A(_09228_),
    .B(_09229_),
    .Y(_09230_));
 sky130_fd_sc_hd__o21ai_2 _23157_ (.A1(_09227_),
    .A2(_09203_),
    .B1(_09230_),
    .Y(_09231_));
 sky130_fd_sc_hd__xnor2_1 _23158_ (.A(_13602_),
    .B(_09231_),
    .Y(\hash.CA1.p1[14] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_646 ();
 sky130_fd_sc_hd__o21ai_0 _23160_ (.A1(_09224_),
    .A2(_09225_),
    .B1(_13598_),
    .Y(_09233_));
 sky130_fd_sc_hd__nand2b_1 _23161_ (.A_N(_13597_),
    .B(_09233_),
    .Y(_09234_));
 sky130_fd_sc_hd__a21oi_1 _23162_ (.A1(_13602_),
    .A2(_09234_),
    .B1(_13601_),
    .Y(_09235_));
 sky130_fd_sc_hd__xnor2_1 _23163_ (.A(_13606_),
    .B(_09235_),
    .Y(\hash.CA1.p1[15] ));
 sky130_fd_sc_hd__inv_1 _23164_ (.A(_13602_),
    .Y(_09236_));
 sky130_fd_sc_hd__o21bai_1 _23165_ (.A1(_09236_),
    .A2(_09231_),
    .B1_N(_13601_),
    .Y(_09237_));
 sky130_fd_sc_hd__a21oi_1 _23166_ (.A1(_13606_),
    .A2(_09237_),
    .B1(_13605_),
    .Y(_09238_));
 sky130_fd_sc_hd__xnor2_1 _23167_ (.A(_13610_),
    .B(_09238_),
    .Y(\hash.CA1.p1[16] ));
 sky130_fd_sc_hd__inv_1 _23168_ (.A(_13606_),
    .Y(_09239_));
 sky130_fd_sc_hd__o21bai_1 _23169_ (.A1(_09239_),
    .A2(_09235_),
    .B1_N(_13605_),
    .Y(_09240_));
 sky130_fd_sc_hd__a21oi_1 _23170_ (.A1(_13610_),
    .A2(_09240_),
    .B1(_13609_),
    .Y(_09241_));
 sky130_fd_sc_hd__xnor2_1 _23171_ (.A(_13614_),
    .B(_09241_),
    .Y(\hash.CA1.p1[17] ));
 sky130_fd_sc_hd__inv_1 _23172_ (.A(_13614_),
    .Y(_09242_));
 sky130_fd_sc_hd__and2_0 _23173_ (.A(_13610_),
    .B(_13605_),
    .X(_09243_));
 sky130_fd_sc_hd__a311oi_1 _23174_ (.A1(_13606_),
    .A2(_09237_),
    .A3(_13610_),
    .B1(_09243_),
    .C1(_13609_),
    .Y(_09244_));
 sky130_fd_sc_hd__o21bai_1 _23175_ (.A1(_09242_),
    .A2(_09244_),
    .B1_N(_13613_),
    .Y(_09245_));
 sky130_fd_sc_hd__xor2_1 _23176_ (.A(_13618_),
    .B(_09245_),
    .X(\hash.CA1.p1[18] ));
 sky130_fd_sc_hd__and3_4 _23177_ (.A(_13610_),
    .B(_13614_),
    .C(_13618_),
    .X(_09246_));
 sky130_fd_sc_hd__a21o_1 _23178_ (.A1(_13606_),
    .A2(_13601_),
    .B1(_13605_),
    .X(_09247_));
 sky130_fd_sc_hd__a21o_1 _23179_ (.A1(_13614_),
    .A2(_13609_),
    .B1(_13613_),
    .X(_09248_));
 sky130_fd_sc_hd__a221oi_4 _23180_ (.A1(_09246_),
    .A2(_09247_),
    .B1(_09248_),
    .B2(_13618_),
    .C1(_13617_),
    .Y(_09249_));
 sky130_fd_sc_hd__clkinv_2 _23181_ (.A(_09249_),
    .Y(_09250_));
 sky130_fd_sc_hd__nand3_1 _23182_ (.A(_13602_),
    .B(_13606_),
    .C(_09246_),
    .Y(_09251_));
 sky130_fd_sc_hd__a21oi_1 _23183_ (.A1(_13598_),
    .A2(_09224_),
    .B1(_13597_),
    .Y(_09252_));
 sky130_fd_sc_hd__nor2_1 _23184_ (.A(_09251_),
    .B(_09252_),
    .Y(_09253_));
 sky130_fd_sc_hd__and3_4 _23185_ (.A(_13602_),
    .B(_13606_),
    .C(_09246_),
    .X(_09254_));
 sky130_fd_sc_hd__nand4_1 _23186_ (.A(_09254_),
    .B(_13590_),
    .C(_13594_),
    .D(_13598_),
    .Y(_09255_));
 sky130_fd_sc_hd__nor3_4 _23187_ (.A(_09207_),
    .B(_09220_),
    .C(_09255_),
    .Y(_09256_));
 sky130_fd_sc_hd__nor3_1 _23188_ (.A(_09250_),
    .B(_09253_),
    .C(_09256_),
    .Y(_09257_));
 sky130_fd_sc_hd__xnor2_1 _23189_ (.A(_13622_),
    .B(_09257_),
    .Y(\hash.CA1.p1[19] ));
 sky130_fd_sc_hd__o21ai_1 _23190_ (.A1(net1111),
    .A2(_09251_),
    .B1(_09249_),
    .Y(_09258_));
 sky130_fd_sc_hd__a21oi_2 _23191_ (.A1(_09258_),
    .A2(_13622_),
    .B1(_13621_),
    .Y(_09259_));
 sky130_fd_sc_hd__xnor2_2 _23192_ (.A(_13626_),
    .B(_09259_),
    .Y(\hash.CA1.p1[20] ));
 sky130_fd_sc_hd__o31ai_4 _23193_ (.A1(_09250_),
    .A2(_09253_),
    .A3(_09256_),
    .B1(_13622_),
    .Y(_09260_));
 sky130_fd_sc_hd__nor2_2 _23194_ (.A(_13621_),
    .B(_13625_),
    .Y(_09261_));
 sky130_fd_sc_hd__nor2_1 _23195_ (.A(_13626_),
    .B(_13625_),
    .Y(_09262_));
 sky130_fd_sc_hd__a21oi_4 _23196_ (.A1(_09261_),
    .A2(_09260_),
    .B1(_09262_),
    .Y(_09263_));
 sky130_fd_sc_hd__xor2_2 _23197_ (.A(_13630_),
    .B(_09263_),
    .X(\hash.CA1.p1[21] ));
 sky130_fd_sc_hd__and3_1 _23198_ (.A(_13622_),
    .B(_13626_),
    .C(_09254_),
    .X(_09264_));
 sky130_fd_sc_hd__o211ai_1 _23199_ (.A1(_09203_),
    .A2(_09227_),
    .B1(_09230_),
    .C1(_09264_),
    .Y(_09265_));
 sky130_fd_sc_hd__and3_4 _23200_ (.A(_13622_),
    .B(_13626_),
    .C(_09250_),
    .X(_09266_));
 sky130_fd_sc_hd__a21oi_2 _23201_ (.A1(_13626_),
    .A2(_13621_),
    .B1(_09266_),
    .Y(_09267_));
 sky130_fd_sc_hd__nand3b_1 _23202_ (.A_N(_13625_),
    .B(_09267_),
    .C(_09265_),
    .Y(_09268_));
 sky130_fd_sc_hd__a21oi_2 _23203_ (.A1(_09268_),
    .A2(_13630_),
    .B1(_13629_),
    .Y(_09269_));
 sky130_fd_sc_hd__xnor2_1 _23204_ (.A(_09269_),
    .B(_13634_),
    .Y(\hash.CA1.p1[22] ));
 sky130_fd_sc_hd__a21o_1 _23205_ (.A1(_09263_),
    .A2(_13630_),
    .B1(_13629_),
    .X(_09270_));
 sky130_fd_sc_hd__a21oi_1 _23206_ (.A1(_13634_),
    .A2(_09270_),
    .B1(_13633_),
    .Y(_09271_));
 sky130_fd_sc_hd__xnor2_1 _23207_ (.A(_09271_),
    .B(_13638_),
    .Y(\hash.CA1.p1[23] ));
 sky130_fd_sc_hd__and3_4 _23208_ (.A(_13630_),
    .B(_13634_),
    .C(_13638_),
    .X(_09272_));
 sky130_fd_sc_hd__a21o_1 _23209_ (.A1(_13634_),
    .A2(_13629_),
    .B1(_13633_),
    .X(_09273_));
 sky130_fd_sc_hd__a21oi_2 _23210_ (.A1(_13638_),
    .A2(_09273_),
    .B1(_13637_),
    .Y(_09274_));
 sky130_fd_sc_hd__a21boi_2 _23211_ (.A1(_09268_),
    .A2(_09272_),
    .B1_N(_09274_),
    .Y(_09275_));
 sky130_fd_sc_hd__xnor2_2 _23212_ (.A(_13642_),
    .B(_09275_),
    .Y(\hash.CA1.p1[24] ));
 sky130_fd_sc_hd__nand2_1 _23213_ (.A(_13642_),
    .B(_13646_),
    .Y(_09276_));
 sky130_fd_sc_hd__nand2_1 _23214_ (.A(_13646_),
    .B(_13641_),
    .Y(_09277_));
 sky130_fd_sc_hd__o21ai_0 _23215_ (.A1(_09274_),
    .A2(_09276_),
    .B1(_09277_),
    .Y(_09278_));
 sky130_fd_sc_hd__a41o_4 _23216_ (.A1(_09263_),
    .A2(_13646_),
    .A3(_13642_),
    .A4(_09272_),
    .B1(_09278_),
    .X(_09279_));
 sky130_fd_sc_hd__nand2_1 _23217_ (.A(_09263_),
    .B(_09272_),
    .Y(_09280_));
 sky130_fd_sc_hd__nand2_1 _23218_ (.A(_09274_),
    .B(_09280_),
    .Y(_09281_));
 sky130_fd_sc_hd__a211oi_2 _23219_ (.A1(_13642_),
    .A2(_09281_),
    .B1(_13641_),
    .C1(_13646_),
    .Y(_09282_));
 sky130_fd_sc_hd__nor2_1 _23220_ (.A(_09279_),
    .B(_09282_),
    .Y(\hash.CA1.p1[25] ));
 sky130_fd_sc_hd__nand4b_1 _23221_ (.A_N(_13625_),
    .B(_09265_),
    .C(_09267_),
    .D(_09274_),
    .Y(_09283_));
 sky130_fd_sc_hd__nand2b_1 _23222_ (.A_N(_09272_),
    .B(_09274_),
    .Y(_09284_));
 sky130_fd_sc_hd__a31o_1 _23223_ (.A1(_13642_),
    .A2(_09283_),
    .A3(_09284_),
    .B1(_13641_),
    .X(_09285_));
 sky130_fd_sc_hd__a21oi_2 _23224_ (.A1(_09285_),
    .A2(_13646_),
    .B1(_13645_),
    .Y(_09286_));
 sky130_fd_sc_hd__xnor2_1 _23225_ (.A(_09286_),
    .B(_13650_),
    .Y(\hash.CA1.p1[26] ));
 sky130_fd_sc_hd__o21a_1 _23226_ (.A1(_13645_),
    .A2(_09279_),
    .B1(_13650_),
    .X(_09287_));
 sky130_fd_sc_hd__nor2_1 _23227_ (.A(_13649_),
    .B(_09287_),
    .Y(_09288_));
 sky130_fd_sc_hd__xnor2_1 _23228_ (.A(_13654_),
    .B(_09288_),
    .Y(\hash.CA1.p1[27] ));
 sky130_fd_sc_hd__a21o_1 _23229_ (.A1(_13638_),
    .A2(_13633_),
    .B1(_13637_),
    .X(_09289_));
 sky130_fd_sc_hd__a21oi_1 _23230_ (.A1(_13642_),
    .A2(_09289_),
    .B1(_13641_),
    .Y(_09290_));
 sky130_fd_sc_hd__nor2b_1 _23231_ (.A(_09290_),
    .B_N(_13646_),
    .Y(_09291_));
 sky130_fd_sc_hd__o21ai_0 _23232_ (.A1(_13645_),
    .A2(_09291_),
    .B1(_13650_),
    .Y(_09292_));
 sky130_fd_sc_hd__nand2b_1 _23233_ (.A_N(_13649_),
    .B(_09292_),
    .Y(_09293_));
 sky130_fd_sc_hd__a21oi_1 _23234_ (.A1(_13654_),
    .A2(_09293_),
    .B1(_13653_),
    .Y(_09294_));
 sky130_fd_sc_hd__nor2_1 _23235_ (.A(_13625_),
    .B(_13629_),
    .Y(_09295_));
 sky130_fd_sc_hd__nand4_1 _23236_ (.A(_09265_),
    .B(_09267_),
    .C(_09294_),
    .D(_09295_),
    .Y(_09296_));
 sky130_fd_sc_hd__nand2_1 _23237_ (.A(_13634_),
    .B(_13638_),
    .Y(_09297_));
 sky130_fd_sc_hd__nand2_1 _23238_ (.A(_13650_),
    .B(_13654_),
    .Y(_09298_));
 sky130_fd_sc_hd__nor2_2 _23239_ (.A(_13630_),
    .B(_13629_),
    .Y(_09299_));
 sky130_fd_sc_hd__o41ai_1 _23240_ (.A1(_09297_),
    .A2(_09276_),
    .A3(_09298_),
    .A4(_09299_),
    .B1(_09294_),
    .Y(_09300_));
 sky130_fd_sc_hd__nand2_1 _23241_ (.A(_09296_),
    .B(_09300_),
    .Y(_09301_));
 sky130_fd_sc_hd__xnor2_2 _23242_ (.A(_13658_),
    .B(_09301_),
    .Y(\hash.CA1.p1[28] ));
 sky130_fd_sc_hd__a21o_4 _23243_ (.A1(_13658_),
    .A2(_13653_),
    .B1(_13657_),
    .X(_09302_));
 sky130_fd_sc_hd__or4_4 _23244_ (.A(_13645_),
    .B(_13649_),
    .C(_09302_),
    .D(_09279_),
    .X(_09303_));
 sky130_fd_sc_hd__a21oi_1 _23245_ (.A1(_13654_),
    .A2(_13658_),
    .B1(_09302_),
    .Y(_09304_));
 sky130_fd_sc_hd__nor3_1 _23246_ (.A(_13650_),
    .B(_13649_),
    .C(_09302_),
    .Y(_09305_));
 sky130_fd_sc_hd__nor2_1 _23247_ (.A(_09304_),
    .B(_09305_),
    .Y(_09306_));
 sky130_fd_sc_hd__nand2_2 _23248_ (.A(_09303_),
    .B(_09306_),
    .Y(_09307_));
 sky130_fd_sc_hd__xnor2_2 _23249_ (.A(_09307_),
    .B(_13662_),
    .Y(\hash.CA1.p1[29] ));
 sky130_fd_sc_hd__xnor2_1 _23250_ (.A(_12882_),
    .B(_13554_),
    .Y(\hash.CA1.p1[2] ));
 sky130_fd_sc_hd__a31o_1 _23251_ (.A1(_13658_),
    .A2(_09296_),
    .A3(_09300_),
    .B1(_13657_),
    .X(_09308_));
 sky130_fd_sc_hd__a21oi_2 _23252_ (.A1(_13662_),
    .A2(_09308_),
    .B1(_13661_),
    .Y(_09309_));
 sky130_fd_sc_hd__xnor2_1 _23253_ (.A(_13666_),
    .B(_09309_),
    .Y(\hash.CA1.p1[30] ));
 sky130_fd_sc_hd__xor2_1 _23254_ (.A(_13241_),
    .B(_06073_),
    .X(_09310_));
 sky130_fd_sc_hd__xnor3_1 _23255_ (.A(\hash.CA2.b_dash[31] ),
    .B(_06248_),
    .C(_06266_),
    .X(_09311_));
 sky130_fd_sc_hd__maj3_1 _23256_ (.A(\hash.CA2.a_dash[31] ),
    .B(net1079),
    .C(_09311_),
    .X(_09312_));
 sky130_fd_sc_hd__xnor2_1 _23257_ (.A(_09310_),
    .B(_09312_),
    .Y(_09313_));
 sky130_fd_sc_hd__nor2_1 _23258_ (.A(net341),
    .B(_09313_),
    .Y(_09314_));
 sky130_fd_sc_hd__inv_1 _23259_ (.A(_13666_),
    .Y(_09315_));
 sky130_fd_sc_hd__a31oi_4 _23260_ (.A1(_09303_),
    .A2(_13662_),
    .A3(_09306_),
    .B1(_13661_),
    .Y(_09316_));
 sky130_fd_sc_hd__o21bai_1 _23261_ (.A1(_09316_),
    .A2(_09315_),
    .B1_N(_13665_),
    .Y(_09317_));
 sky130_fd_sc_hd__xor2_1 _23262_ (.A(_06156_),
    .B(_09317_),
    .X(_09318_));
 sky130_fd_sc_hd__xnor2_1 _23263_ (.A(_09314_),
    .B(_09318_),
    .Y(\hash.CA1.p1[31] ));
 sky130_fd_sc_hd__xnor2_1 _23264_ (.A(_13558_),
    .B(_09210_),
    .Y(\hash.CA1.p1[3] ));
 sky130_fd_sc_hd__nand2_1 _23265_ (.A(_09194_),
    .B(_09196_),
    .Y(_09319_));
 sky130_fd_sc_hd__nor2_1 _23266_ (.A(_13562_),
    .B(_09319_),
    .Y(_09320_));
 sky130_fd_sc_hd__nor2_2 _23267_ (.A(_09197_),
    .B(_09320_),
    .Y(\hash.CA1.p1[4] ));
 sky130_fd_sc_hd__o21ai_0 _23268_ (.A1(_09208_),
    .A2(_09210_),
    .B1(_09194_),
    .Y(_09321_));
 sky130_fd_sc_hd__a21oi_1 _23269_ (.A1(_13562_),
    .A2(_09321_),
    .B1(_13561_),
    .Y(_09322_));
 sky130_fd_sc_hd__xnor2_1 _23270_ (.A(_13566_),
    .B(_09322_),
    .Y(\hash.CA1.p1[5] ));
 sky130_fd_sc_hd__nand2_1 _23271_ (.A(_09193_),
    .B(_09198_),
    .Y(_09323_));
 sky130_fd_sc_hd__nor2_1 _23272_ (.A(_13570_),
    .B(_09323_),
    .Y(_09324_));
 sky130_fd_sc_hd__nor2_2 _23273_ (.A(_09199_),
    .B(_09324_),
    .Y(\hash.CA1.p1[6] ));
 sky130_fd_sc_hd__a31oi_1 _23274_ (.A1(_13570_),
    .A2(_09212_),
    .A3(_09214_),
    .B1(_13569_),
    .Y(_09325_));
 sky130_fd_sc_hd__xnor2_1 _23275_ (.A(_13574_),
    .B(_09325_),
    .Y(\hash.CA1.p1[7] ));
 sky130_fd_sc_hd__nand2_1 _23276_ (.A(_09192_),
    .B(_09200_),
    .Y(_09326_));
 sky130_fd_sc_hd__nor2_1 _23277_ (.A(_13578_),
    .B(_09326_),
    .Y(_09327_));
 sky130_fd_sc_hd__nor2_4 _23278_ (.A(_09201_),
    .B(_09327_),
    .Y(\hash.CA1.p1[8] ));
 sky130_fd_sc_hd__nand2b_2 _23279_ (.A_N(_09216_),
    .B(_09219_),
    .Y(_09328_));
 sky130_fd_sc_hd__xor2_2 _23280_ (.A(_13582_),
    .B(_09328_),
    .X(\hash.CA1.p1[9] ));
 sky130_fd_sc_hd__inv_1 _23281_ (.A(_14155_),
    .Y(_09329_));
 sky130_fd_sc_hd__inv_1 _23282_ (.A(_14147_),
    .Y(_09330_));
 sky130_fd_sc_hd__a21o_1 _23283_ (.A1(_14207_),
    .A2(_14131_),
    .B1(_14130_),
    .X(_09331_));
 sky130_fd_sc_hd__a21o_4 _23284_ (.A1(_14135_),
    .A2(_09331_),
    .B1(_14134_),
    .X(_09332_));
 sky130_fd_sc_hd__a21oi_1 _23285_ (.A1(_14139_),
    .A2(_09332_),
    .B1(_14138_),
    .Y(_09333_));
 sky130_fd_sc_hd__nor2b_1 _23286_ (.A(_09333_),
    .B_N(_14143_),
    .Y(_09334_));
 sky130_fd_sc_hd__nor2_2 _23287_ (.A(_14142_),
    .B(_09334_),
    .Y(_09335_));
 sky130_fd_sc_hd__o21bai_1 _23288_ (.A1(_09330_),
    .A2(_09335_),
    .B1_N(_14146_),
    .Y(_09336_));
 sky130_fd_sc_hd__a21oi_2 _23289_ (.A1(_14151_),
    .A2(_09336_),
    .B1(_14150_),
    .Y(_09337_));
 sky130_fd_sc_hd__o21bai_1 _23290_ (.A1(_09329_),
    .A2(_09337_),
    .B1_N(_14154_),
    .Y(_09338_));
 sky130_fd_sc_hd__a21oi_1 _23291_ (.A1(_14158_),
    .A2(_09338_),
    .B1(_14157_),
    .Y(_09339_));
 sky130_fd_sc_hd__xnor2_1 _23292_ (.A(_14160_),
    .B(_09339_),
    .Y(\hash.CA1.p2[10] ));
 sky130_fd_sc_hd__a21o_1 _23293_ (.A1(_14158_),
    .A2(_14154_),
    .B1(_14157_),
    .X(_09340_));
 sky130_fd_sc_hd__a21o_4 _23294_ (.A1(_14160_),
    .A2(_09340_),
    .B1(_14159_),
    .X(_09341_));
 sky130_fd_sc_hd__nor2b_1 _23295_ (.A(_12885_),
    .B_N(_14135_),
    .Y(_09342_));
 sky130_fd_sc_hd__o21a_1 _23296_ (.A1(_14134_),
    .A2(_09342_),
    .B1(_14139_),
    .X(_09343_));
 sky130_fd_sc_hd__o21ai_2 _23297_ (.A1(_14138_),
    .A2(_09343_),
    .B1(_14143_),
    .Y(_09344_));
 sky130_fd_sc_hd__nor3_1 _23298_ (.A(_14142_),
    .B(_14146_),
    .C(_14150_),
    .Y(_09345_));
 sky130_fd_sc_hd__inv_1 _23299_ (.A(_14151_),
    .Y(_09346_));
 sky130_fd_sc_hd__nor2_1 _23300_ (.A(_14147_),
    .B(_14146_),
    .Y(_09347_));
 sky130_fd_sc_hd__nor2_1 _23301_ (.A(_09346_),
    .B(_09347_),
    .Y(_09348_));
 sky130_fd_sc_hd__and3_4 _23302_ (.A(_14160_),
    .B(_14155_),
    .C(_14158_),
    .X(_09349_));
 sky130_fd_sc_hd__o21ai_2 _23303_ (.A1(_14150_),
    .A2(_09348_),
    .B1(_09349_),
    .Y(_09350_));
 sky130_fd_sc_hd__a21oi_2 _23304_ (.A1(_09344_),
    .A2(_09345_),
    .B1(_09350_),
    .Y(_09351_));
 sky130_fd_sc_hd__nor2_1 _23305_ (.A(_09341_),
    .B(_09351_),
    .Y(_09352_));
 sky130_fd_sc_hd__xnor2_1 _23306_ (.A(_14162_),
    .B(_09352_),
    .Y(\hash.CA1.p2[11] ));
 sky130_fd_sc_hd__a211oi_1 _23307_ (.A1(_14139_),
    .A2(_09332_),
    .B1(_14142_),
    .C1(_14138_),
    .Y(_09353_));
 sky130_fd_sc_hd__o2111ai_2 _23308_ (.A1(_14143_),
    .A2(_14142_),
    .B1(_14151_),
    .C1(_14147_),
    .D1(_09349_),
    .Y(_09354_));
 sky130_fd_sc_hd__a21o_1 _23309_ (.A1(_14151_),
    .A2(_14146_),
    .B1(_14150_),
    .X(_09355_));
 sky130_fd_sc_hd__a21oi_2 _23310_ (.A1(_09349_),
    .A2(_09355_),
    .B1(_09341_),
    .Y(_09356_));
 sky130_fd_sc_hd__o21ai_2 _23311_ (.A1(_09353_),
    .A2(_09354_),
    .B1(_09356_),
    .Y(_09357_));
 sky130_fd_sc_hd__a21oi_1 _23312_ (.A1(_14162_),
    .A2(_09357_),
    .B1(_14161_),
    .Y(_09358_));
 sky130_fd_sc_hd__xnor2_2 _23313_ (.A(_14164_),
    .B(_09358_),
    .Y(\hash.CA1.p2[12] ));
 sky130_fd_sc_hd__inv_1 _23314_ (.A(_14161_),
    .Y(_09359_));
 sky130_fd_sc_hd__o21ai_4 _23315_ (.A1(_09341_),
    .A2(_09351_),
    .B1(_14162_),
    .Y(_09360_));
 sky130_fd_sc_hd__nand2_1 _23316_ (.A(_09359_),
    .B(_09360_),
    .Y(_09361_));
 sky130_fd_sc_hd__a21o_4 _23317_ (.A1(_14164_),
    .A2(_09361_),
    .B1(_14163_),
    .X(_09362_));
 sky130_fd_sc_hd__xor2_2 _23318_ (.A(_14166_),
    .B(_09362_),
    .X(\hash.CA1.p2[13] ));
 sky130_fd_sc_hd__nor3_2 _23319_ (.A(_14161_),
    .B(_14163_),
    .C(_09357_),
    .Y(_09363_));
 sky130_fd_sc_hd__o21a_1 _23320_ (.A1(_14162_),
    .A2(_14161_),
    .B1(_14164_),
    .X(_09364_));
 sky130_fd_sc_hd__nor2_1 _23321_ (.A(_14163_),
    .B(_09364_),
    .Y(_09365_));
 sky130_fd_sc_hd__nor2_1 _23322_ (.A(_09363_),
    .B(_09365_),
    .Y(_09366_));
 sky130_fd_sc_hd__a21oi_1 _23323_ (.A1(_14166_),
    .A2(_09366_),
    .B1(_14165_),
    .Y(_09367_));
 sky130_fd_sc_hd__xnor2_2 _23324_ (.A(_14168_),
    .B(_09367_),
    .Y(\hash.CA1.p2[14] ));
 sky130_fd_sc_hd__a21o_1 _23325_ (.A1(_14166_),
    .A2(_09362_),
    .B1(_14165_),
    .X(_09368_));
 sky130_fd_sc_hd__a21oi_1 _23326_ (.A1(_14168_),
    .A2(_09368_),
    .B1(_14167_),
    .Y(_09369_));
 sky130_fd_sc_hd__xnor2_1 _23327_ (.A(_14170_),
    .B(_09369_),
    .Y(\hash.CA1.p2[15] ));
 sky130_fd_sc_hd__nand3_1 _23328_ (.A(_14166_),
    .B(_14168_),
    .C(_14170_),
    .Y(_09370_));
 sky130_fd_sc_hd__or3_4 _23329_ (.A(_09363_),
    .B(_09365_),
    .C(_09370_),
    .X(_09371_));
 sky130_fd_sc_hd__a21o_1 _23330_ (.A1(_14168_),
    .A2(_14165_),
    .B1(_14167_),
    .X(_09372_));
 sky130_fd_sc_hd__a21oi_4 _23331_ (.A1(_14170_),
    .A2(_09372_),
    .B1(_14169_),
    .Y(_09373_));
 sky130_fd_sc_hd__nand2_1 _23332_ (.A(_09371_),
    .B(_09373_),
    .Y(_09374_));
 sky130_fd_sc_hd__xor2_1 _23333_ (.A(_14172_),
    .B(_09374_),
    .X(\hash.CA1.p2[16] ));
 sky130_fd_sc_hd__nand4_1 _23334_ (.A(_14164_),
    .B(_14166_),
    .C(_14168_),
    .D(_14170_),
    .Y(_09375_));
 sky130_fd_sc_hd__a21oi_2 _23335_ (.A1(_09359_),
    .A2(_09360_),
    .B1(_09375_),
    .Y(_09376_));
 sky130_fd_sc_hd__nand4_1 _23336_ (.A(_14166_),
    .B(_14168_),
    .C(_14170_),
    .D(_14163_),
    .Y(_09377_));
 sky130_fd_sc_hd__nand2_1 _23337_ (.A(_09373_),
    .B(_09377_),
    .Y(_09378_));
 sky130_fd_sc_hd__o21a_1 _23338_ (.A1(_09376_),
    .A2(_09378_),
    .B1(_14172_),
    .X(_09379_));
 sky130_fd_sc_hd__nor2_1 _23339_ (.A(_14171_),
    .B(_09379_),
    .Y(_09380_));
 sky130_fd_sc_hd__xnor2_1 _23340_ (.A(_14174_),
    .B(_09380_),
    .Y(\hash.CA1.p2[17] ));
 sky130_fd_sc_hd__nor2_1 _23341_ (.A(_14171_),
    .B(_14173_),
    .Y(_09381_));
 sky130_fd_sc_hd__o21a_1 _23342_ (.A1(_14172_),
    .A2(_14171_),
    .B1(_14174_),
    .X(_09382_));
 sky130_fd_sc_hd__nor2_1 _23343_ (.A(_14173_),
    .B(_09382_),
    .Y(_09383_));
 sky130_fd_sc_hd__a31oi_4 _23344_ (.A1(_09371_),
    .A2(_09373_),
    .A3(_09381_),
    .B1(_09383_),
    .Y(_09384_));
 sky130_fd_sc_hd__xor2_1 _23345_ (.A(_14176_),
    .B(_09384_),
    .X(\hash.CA1.p2[18] ));
 sky130_fd_sc_hd__o2111ai_2 _23346_ (.A1(_09376_),
    .A2(_09378_),
    .B1(_14172_),
    .C1(_14174_),
    .D1(_14176_),
    .Y(_09385_));
 sky130_fd_sc_hd__and3_1 _23347_ (.A(_14174_),
    .B(_14176_),
    .C(_14171_),
    .X(_09386_));
 sky130_fd_sc_hd__a21oi_1 _23348_ (.A1(_14176_),
    .A2(_14173_),
    .B1(_09386_),
    .Y(_09387_));
 sky130_fd_sc_hd__nand3b_1 _23349_ (.A_N(_14175_),
    .B(_09385_),
    .C(_09387_),
    .Y(_09388_));
 sky130_fd_sc_hd__xor2_1 _23350_ (.A(_14178_),
    .B(_09388_),
    .X(\hash.CA1.p2[19] ));
 sky130_fd_sc_hd__nand2_1 _23351_ (.A(_14180_),
    .B(_14177_),
    .Y(_09389_));
 sky130_fd_sc_hd__nand3_1 _23352_ (.A(_14178_),
    .B(_14180_),
    .C(_14175_),
    .Y(_09390_));
 sky130_fd_sc_hd__nand2_1 _23353_ (.A(_09389_),
    .B(_09390_),
    .Y(_09391_));
 sky130_fd_sc_hd__a41o_4 _23354_ (.A1(_09384_),
    .A2(_14178_),
    .A3(_14180_),
    .A4(_14176_),
    .B1(_09391_),
    .X(_09392_));
 sky130_fd_sc_hd__a21o_1 _23355_ (.A1(_14176_),
    .A2(_09384_),
    .B1(_14175_),
    .X(_09393_));
 sky130_fd_sc_hd__a211oi_1 _23356_ (.A1(_14178_),
    .A2(_09393_),
    .B1(_14177_),
    .C1(_14180_),
    .Y(_09394_));
 sky130_fd_sc_hd__nor2_1 _23357_ (.A(_09392_),
    .B(_09394_),
    .Y(\hash.CA1.p2[20] ));
 sky130_fd_sc_hd__nor3_1 _23358_ (.A(_14175_),
    .B(_14177_),
    .C(_14179_),
    .Y(_09395_));
 sky130_fd_sc_hd__or2_0 _23359_ (.A(_14178_),
    .B(_14177_),
    .X(_09396_));
 sky130_fd_sc_hd__a21oi_1 _23360_ (.A1(_14180_),
    .A2(_09396_),
    .B1(_14179_),
    .Y(_09397_));
 sky130_fd_sc_hd__a31oi_2 _23361_ (.A1(_09395_),
    .A2(_09385_),
    .A3(_09387_),
    .B1(_09397_),
    .Y(_09398_));
 sky130_fd_sc_hd__and2_4 _23362_ (.A(_14182_),
    .B(_09398_),
    .X(_09399_));
 sky130_fd_sc_hd__nor2_1 _23363_ (.A(_14182_),
    .B(_09398_),
    .Y(_09400_));
 sky130_fd_sc_hd__nor2_1 _23364_ (.A(_09399_),
    .B(_09400_),
    .Y(\hash.CA1.p2[21] ));
 sky130_fd_sc_hd__o21a_1 _23365_ (.A1(_14179_),
    .A2(_09392_),
    .B1(_14182_),
    .X(_09401_));
 sky130_fd_sc_hd__nor2_1 _23366_ (.A(_14181_),
    .B(_09401_),
    .Y(_09402_));
 sky130_fd_sc_hd__xnor2_1 _23367_ (.A(_14184_),
    .B(_09402_),
    .Y(\hash.CA1.p2[22] ));
 sky130_fd_sc_hd__inv_2 _23368_ (.A(_14183_),
    .Y(_09403_));
 sky130_fd_sc_hd__o21ai_4 _23369_ (.A1(_14181_),
    .A2(_09399_),
    .B1(_14184_),
    .Y(_09404_));
 sky130_fd_sc_hd__clkinv_1 _23370_ (.A(_14186_),
    .Y(_09405_));
 sky130_fd_sc_hd__a21oi_4 _23371_ (.A1(_09403_),
    .A2(_09404_),
    .B1(_09405_),
    .Y(_09406_));
 sky130_fd_sc_hd__and3_1 _23372_ (.A(_09405_),
    .B(_09403_),
    .C(_09404_),
    .X(_09407_));
 sky130_fd_sc_hd__nor2_1 _23373_ (.A(_09407_),
    .B(_09406_),
    .Y(\hash.CA1.p2[23] ));
 sky130_fd_sc_hd__inv_1 _23374_ (.A(_14184_),
    .Y(_09408_));
 sky130_fd_sc_hd__nor2_1 _23375_ (.A(_14182_),
    .B(_14181_),
    .Y(_09409_));
 sky130_fd_sc_hd__o21ai_0 _23376_ (.A1(_09408_),
    .A2(_09409_),
    .B1(_09403_),
    .Y(_09410_));
 sky130_fd_sc_hd__o41ai_4 _23377_ (.A1(_14179_),
    .A2(_14181_),
    .A3(_14183_),
    .A4(_09392_),
    .B1(_09410_),
    .Y(_09411_));
 sky130_fd_sc_hd__o21bai_1 _23378_ (.A1(_09405_),
    .A2(_09411_),
    .B1_N(_14185_),
    .Y(_09412_));
 sky130_fd_sc_hd__xor2_1 _23379_ (.A(_14188_),
    .B(_09412_),
    .X(\hash.CA1.p2[24] ));
 sky130_fd_sc_hd__o21a_1 _23380_ (.A1(_14185_),
    .A2(_09406_),
    .B1(_14188_),
    .X(_09413_));
 sky130_fd_sc_hd__nor2_1 _23381_ (.A(_14187_),
    .B(_09413_),
    .Y(_09414_));
 sky130_fd_sc_hd__xnor2_1 _23382_ (.A(_14190_),
    .B(_09414_),
    .Y(\hash.CA1.p2[25] ));
 sky130_fd_sc_hd__nand3_1 _23383_ (.A(_14186_),
    .B(_14188_),
    .C(_14190_),
    .Y(_09415_));
 sky130_fd_sc_hd__a21oi_4 _23384_ (.A1(_14188_),
    .A2(_14185_),
    .B1(_14187_),
    .Y(_09416_));
 sky130_fd_sc_hd__inv_1 _23385_ (.A(_14190_),
    .Y(_09417_));
 sky130_fd_sc_hd__o22ai_2 _23386_ (.A1(_09411_),
    .A2(_09415_),
    .B1(_09416_),
    .B2(_09417_),
    .Y(_09418_));
 sky130_fd_sc_hd__nor2_2 _23387_ (.A(_09418_),
    .B(_14189_),
    .Y(_09419_));
 sky130_fd_sc_hd__xnor2_1 _23388_ (.A(_14192_),
    .B(_09419_),
    .Y(\hash.CA1.p2[26] ));
 sky130_fd_sc_hd__nor2_1 _23389_ (.A(_14188_),
    .B(_14187_),
    .Y(_09420_));
 sky130_fd_sc_hd__o21bai_1 _23390_ (.A1(_09417_),
    .A2(_09420_),
    .B1_N(_14189_),
    .Y(_09421_));
 sky130_fd_sc_hd__o41a_1 _23391_ (.A1(_14185_),
    .A2(_14187_),
    .A3(_14189_),
    .A4(_09406_),
    .B1(_09421_),
    .X(_09422_));
 sky130_fd_sc_hd__a21oi_2 _23392_ (.A1(_09422_),
    .A2(_14192_),
    .B1(_14191_),
    .Y(_09423_));
 sky130_fd_sc_hd__xnor2_1 _23393_ (.A(_14194_),
    .B(_09423_),
    .Y(\hash.CA1.p2[27] ));
 sky130_fd_sc_hd__nor3_1 _23394_ (.A(_14192_),
    .B(_14191_),
    .C(_14193_),
    .Y(_09424_));
 sky130_fd_sc_hd__nor2_1 _23395_ (.A(_14194_),
    .B(_14193_),
    .Y(_09425_));
 sky130_fd_sc_hd__nor2_1 _23396_ (.A(_09424_),
    .B(_09425_),
    .Y(_09426_));
 sky130_fd_sc_hd__o41ai_2 _23397_ (.A1(_14189_),
    .A2(_14191_),
    .A3(_14193_),
    .A4(_09418_),
    .B1(_09426_),
    .Y(_09427_));
 sky130_fd_sc_hd__xnor2_1 _23398_ (.A(_14196_),
    .B(_09427_),
    .Y(\hash.CA1.p2[28] ));
 sky130_fd_sc_hd__clkinv_1 _23399_ (.A(_14196_),
    .Y(_09428_));
 sky130_fd_sc_hd__a21oi_1 _23400_ (.A1(_14194_),
    .A2(_14191_),
    .B1(_14193_),
    .Y(_09429_));
 sky130_fd_sc_hd__o21bai_1 _23401_ (.A1(_09428_),
    .A2(_09429_),
    .B1_N(_14195_),
    .Y(_09430_));
 sky130_fd_sc_hd__a41o_1 _23402_ (.A1(_14194_),
    .A2(_09422_),
    .A3(_14196_),
    .A4(_14192_),
    .B1(_09430_),
    .X(_09431_));
 sky130_fd_sc_hd__xor2_1 _23403_ (.A(_14198_),
    .B(_09431_),
    .X(\hash.CA1.p2[29] ));
 sky130_fd_sc_hd__o21bai_1 _23404_ (.A1(_09427_),
    .A2(_09428_),
    .B1_N(_14195_),
    .Y(_09432_));
 sky130_fd_sc_hd__a21oi_2 _23405_ (.A1(_14198_),
    .A2(_09432_),
    .B1(_14197_),
    .Y(_09433_));
 sky130_fd_sc_hd__xnor2_1 _23406_ (.A(_14201_),
    .B(_09433_),
    .Y(\hash.CA1.p2[30] ));
 sky130_fd_sc_hd__xnor2_1 _23407_ (.A(\hash.CA2.f_dash[31] ),
    .B(_08094_),
    .Y(_09434_));
 sky130_fd_sc_hd__nor2_1 _23408_ (.A(net534),
    .B(_09434_),
    .Y(_09435_));
 sky130_fd_sc_hd__xor2_2 _23409_ (.A(\hash.CA1.w_i1[31] ),
    .B(\hash.CA1.k_i1[31] ),
    .X(_09436_));
 sky130_fd_sc_hd__xnor2_1 _23410_ (.A(_09435_),
    .B(_09436_),
    .Y(_09437_));
 sky130_fd_sc_hd__xnor2_1 _23411_ (.A(\hash.CA1.S1.X[10] ),
    .B(_09437_),
    .Y(_09438_));
 sky130_fd_sc_hd__xnor2_1 _23412_ (.A(_06673_),
    .B(_09438_),
    .Y(_09439_));
 sky130_fd_sc_hd__nand2_1 _23413_ (.A(_14115_),
    .B(_14124_),
    .Y(_09440_));
 sky130_fd_sc_hd__a21oi_1 _23414_ (.A1(_14124_),
    .A2(_14114_),
    .B1(_14123_),
    .Y(_09441_));
 sky130_fd_sc_hd__o21ai_0 _23415_ (.A1(_07134_),
    .A2(_09440_),
    .B1(_09441_),
    .Y(_09442_));
 sky130_fd_sc_hd__xnor2_1 _23416_ (.A(_09439_),
    .B(_09442_),
    .Y(_09443_));
 sky130_fd_sc_hd__nor2b_1 _23417_ (.A(_07108_),
    .B_N(_14120_),
    .Y(_09444_));
 sky130_fd_sc_hd__a311oi_1 _23418_ (.A1(_14111_),
    .A2(_14120_),
    .A3(_08101_),
    .B1(_09444_),
    .C1(_14119_),
    .Y(_09445_));
 sky130_fd_sc_hd__xnor2_1 _23419_ (.A(_09443_),
    .B(_09445_),
    .Y(_09446_));
 sky130_fd_sc_hd__nor2b_4 _23420_ (.A(net534),
    .B_N(\hash.CA2.S1.X[31] ),
    .Y(_09447_));
 sky130_fd_sc_hd__mux2i_4 _23421_ (.A0(_09447_),
    .A1(_06418_),
    .S(net1043),
    .Y(_09448_));
 sky130_fd_sc_hd__xnor2_2 _23422_ (.A(_09446_),
    .B(_09448_),
    .Y(_09449_));
 sky130_fd_sc_hd__xor2_1 _23423_ (.A(_12877_),
    .B(_12873_),
    .X(_09450_));
 sky130_fd_sc_hd__nor2_2 _23424_ (.A(net534),
    .B(\hash.CA2.b_dash[31] ),
    .Y(_09451_));
 sky130_fd_sc_hd__xnor2_1 _23425_ (.A(_09450_),
    .B(_09451_),
    .Y(_09452_));
 sky130_fd_sc_hd__nand3_1 _23426_ (.A(_14192_),
    .B(_14194_),
    .C(_14196_),
    .Y(_09453_));
 sky130_fd_sc_hd__nand4_1 _23427_ (.A(_14188_),
    .B(_14190_),
    .C(_14198_),
    .D(_14201_),
    .Y(_09454_));
 sky130_fd_sc_hd__nor2_1 _23428_ (.A(_09453_),
    .B(_09454_),
    .Y(_09455_));
 sky130_fd_sc_hd__nor2_1 _23429_ (.A(_09417_),
    .B(_09416_),
    .Y(_09456_));
 sky130_fd_sc_hd__o21ai_0 _23430_ (.A1(_14189_),
    .A2(_09456_),
    .B1(_14192_),
    .Y(_09457_));
 sky130_fd_sc_hd__nand2b_1 _23431_ (.A_N(_14191_),
    .B(_09457_),
    .Y(_09458_));
 sky130_fd_sc_hd__a21oi_1 _23432_ (.A1(_14194_),
    .A2(_09458_),
    .B1(_14193_),
    .Y(_09459_));
 sky130_fd_sc_hd__o21bai_1 _23433_ (.A1(_09428_),
    .A2(_09459_),
    .B1_N(_14195_),
    .Y(_09460_));
 sky130_fd_sc_hd__a21oi_1 _23434_ (.A1(_14198_),
    .A2(_09460_),
    .B1(_14197_),
    .Y(_09461_));
 sky130_fd_sc_hd__nor2b_1 _23435_ (.A(_09461_),
    .B_N(_14201_),
    .Y(_09462_));
 sky130_fd_sc_hd__a211oi_2 _23436_ (.A1(_09406_),
    .A2(_09455_),
    .B1(_14200_),
    .C1(_09462_),
    .Y(_09463_));
 sky130_fd_sc_hd__xnor2_1 _23437_ (.A(_09452_),
    .B(_09463_),
    .Y(_09464_));
 sky130_fd_sc_hd__xnor2_1 _23438_ (.A(_09449_),
    .B(_09464_),
    .Y(\hash.CA1.p2[31] ));
 sky130_fd_sc_hd__xnor2_1 _23439_ (.A(_12885_),
    .B(_14135_),
    .Y(\hash.CA1.p2[3] ));
 sky130_fd_sc_hd__xor2_1 _23440_ (.A(_14139_),
    .B(_09332_),
    .X(\hash.CA1.p2[4] ));
 sky130_fd_sc_hd__nor2_1 _23441_ (.A(_14138_),
    .B(_09343_),
    .Y(_09465_));
 sky130_fd_sc_hd__xnor2_1 _23442_ (.A(_14143_),
    .B(_09465_),
    .Y(\hash.CA1.p2[5] ));
 sky130_fd_sc_hd__xnor2_2 _23443_ (.A(_14147_),
    .B(_09335_),
    .Y(\hash.CA1.p2[6] ));
 sky130_fd_sc_hd__nand2b_1 _23444_ (.A_N(_14142_),
    .B(_09344_),
    .Y(_09466_));
 sky130_fd_sc_hd__a21oi_2 _23445_ (.A1(_14147_),
    .A2(_09466_),
    .B1(_14146_),
    .Y(_09467_));
 sky130_fd_sc_hd__xnor2_2 _23446_ (.A(_14151_),
    .B(_09467_),
    .Y(\hash.CA1.p2[7] ));
 sky130_fd_sc_hd__xnor2_2 _23447_ (.A(_14155_),
    .B(_09337_),
    .Y(\hash.CA1.p2[8] ));
 sky130_fd_sc_hd__o21bai_1 _23448_ (.A1(_09346_),
    .A2(_09467_),
    .B1_N(_14150_),
    .Y(_09468_));
 sky130_fd_sc_hd__a21oi_1 _23449_ (.A1(_14155_),
    .A2(_09468_),
    .B1(_14154_),
    .Y(_09469_));
 sky130_fd_sc_hd__xnor2_2 _23450_ (.A(_14158_),
    .B(_09469_),
    .Y(\hash.CA1.p2[9] ));
 sky130_fd_sc_hd__clkinvlp_4 _23451_ (.A(_13918_),
    .Y(_09470_));
 sky130_fd_sc_hd__inv_1 _23452_ (.A(_13893_),
    .Y(_09471_));
 sky130_fd_sc_hd__a21o_4 _23453_ (.A1(_14208_),
    .A2(_13874_),
    .B1(_13873_),
    .X(_09472_));
 sky130_fd_sc_hd__a21oi_4 _23454_ (.A1(_13883_),
    .A2(_09472_),
    .B1(_13882_),
    .Y(_09473_));
 sky130_fd_sc_hd__inv_2 _23455_ (.A(_13892_),
    .Y(_09474_));
 sky130_fd_sc_hd__o21ai_0 _23456_ (.A1(_09471_),
    .A2(_09473_),
    .B1(_09474_),
    .Y(_09475_));
 sky130_fd_sc_hd__a21o_4 _23457_ (.A1(_13902_),
    .A2(_09475_),
    .B1(_13901_),
    .X(_09476_));
 sky130_fd_sc_hd__a21oi_4 _23458_ (.A1(_13910_),
    .A2(_09476_),
    .B1(_13909_),
    .Y(_09477_));
 sky130_fd_sc_hd__nor2_1 _23459_ (.A(_09470_),
    .B(_09477_),
    .Y(_09478_));
 sky130_fd_sc_hd__o21ai_0 _23460_ (.A1(_13917_),
    .A2(_09478_),
    .B1(_13927_),
    .Y(_09479_));
 sky130_fd_sc_hd__nand2b_1 _23461_ (.A_N(_13926_),
    .B(_09479_),
    .Y(_09480_));
 sky130_fd_sc_hd__a21oi_2 _23462_ (.A1(_13936_),
    .A2(_09480_),
    .B1(_13935_),
    .Y(_09481_));
 sky130_fd_sc_hd__xnor2_4 _23463_ (.A(_13945_),
    .B(_09481_),
    .Y(\hash.CA1.p3[10] ));
 sky130_fd_sc_hd__nor2b_1 _23464_ (.A(_12892_),
    .B_N(_13883_),
    .Y(_09482_));
 sky130_fd_sc_hd__o21ai_2 _23465_ (.A1(_13882_),
    .A2(_09482_),
    .B1(_13893_),
    .Y(_09483_));
 sky130_fd_sc_hd__a21boi_4 _23466_ (.A1(_09474_),
    .A2(_09483_),
    .B1_N(_13902_),
    .Y(_09484_));
 sky130_fd_sc_hd__nor2_2 _23467_ (.A(_13901_),
    .B(_09484_),
    .Y(_09485_));
 sky130_fd_sc_hd__nand2_1 _23468_ (.A(_13910_),
    .B(_13918_),
    .Y(_09486_));
 sky130_fd_sc_hd__a21oi_1 _23469_ (.A1(_13918_),
    .A2(_13909_),
    .B1(_13917_),
    .Y(_09487_));
 sky130_fd_sc_hd__o21ai_2 _23470_ (.A1(_09485_),
    .A2(_09486_),
    .B1(_09487_),
    .Y(_09488_));
 sky130_fd_sc_hd__and2_4 _23471_ (.A(_13927_),
    .B(_09488_),
    .X(_09489_));
 sky130_fd_sc_hd__o21a_4 _23472_ (.A1(_13926_),
    .A2(_09489_),
    .B1(_13936_),
    .X(_09490_));
 sky130_fd_sc_hd__o21a_4 _23473_ (.A1(_13935_),
    .A2(_09490_),
    .B1(_13945_),
    .X(_09491_));
 sky130_fd_sc_hd__nor2_4 _23474_ (.A(_13944_),
    .B(_09491_),
    .Y(_09492_));
 sky130_fd_sc_hd__xnor2_4 _23475_ (.A(_13955_),
    .B(_09492_),
    .Y(\hash.CA1.p3[11] ));
 sky130_fd_sc_hd__nand4_1 _23476_ (.A(_13945_),
    .B(_13955_),
    .C(_13927_),
    .D(_13936_),
    .Y(_09493_));
 sky130_fd_sc_hd__inv_1 _23477_ (.A(_13955_),
    .Y(_09494_));
 sky130_fd_sc_hd__a21o_1 _23478_ (.A1(_13936_),
    .A2(_13926_),
    .B1(_13935_),
    .X(_09495_));
 sky130_fd_sc_hd__a21oi_2 _23479_ (.A1(_09495_),
    .A2(_13945_),
    .B1(_13944_),
    .Y(_09496_));
 sky130_fd_sc_hd__nor2_2 _23480_ (.A(_09494_),
    .B(_09496_),
    .Y(_09497_));
 sky130_fd_sc_hd__inv_1 _23481_ (.A(_13917_),
    .Y(_09498_));
 sky130_fd_sc_hd__nor2_1 _23482_ (.A(_09493_),
    .B(_09498_),
    .Y(_09499_));
 sky130_fd_sc_hd__nor2_2 _23483_ (.A(_09499_),
    .B(_09497_),
    .Y(_09500_));
 sky130_fd_sc_hd__o31ai_4 _23484_ (.A1(_09470_),
    .A2(_09477_),
    .A3(_09493_),
    .B1(_09500_),
    .Y(_09501_));
 sky130_fd_sc_hd__nor2_2 _23485_ (.A(_13954_),
    .B(_09501_),
    .Y(_09502_));
 sky130_fd_sc_hd__xnor2_4 _23486_ (.A(_13964_),
    .B(_09502_),
    .Y(\hash.CA1.p3[12] ));
 sky130_fd_sc_hd__o21bai_1 _23487_ (.A1(_09494_),
    .A2(_09492_),
    .B1_N(_13954_),
    .Y(_09503_));
 sky130_fd_sc_hd__a21oi_2 _23488_ (.A1(_13964_),
    .A2(_09503_),
    .B1(_13963_),
    .Y(_09504_));
 sky130_fd_sc_hd__xnor2_4 _23489_ (.A(_13972_),
    .B(_09504_),
    .Y(\hash.CA1.p3[13] ));
 sky130_fd_sc_hd__o21ai_0 _23490_ (.A1(_13954_),
    .A2(_09501_),
    .B1(_13964_),
    .Y(_09505_));
 sky130_fd_sc_hd__nand2b_1 _23491_ (.A_N(_13963_),
    .B(_09505_),
    .Y(_09506_));
 sky130_fd_sc_hd__a21oi_1 _23492_ (.A1(_13972_),
    .A2(_09506_),
    .B1(_13971_),
    .Y(_09507_));
 sky130_fd_sc_hd__xnor2_1 _23493_ (.A(_13981_),
    .B(_09507_),
    .Y(\hash.CA1.p3[14] ));
 sky130_fd_sc_hd__o211ai_1 _23494_ (.A1(_13963_),
    .A2(_13964_),
    .B1(_13981_),
    .C1(_13972_),
    .Y(_09508_));
 sky130_fd_sc_hd__nor3_2 _23495_ (.A(_13954_),
    .B(_09497_),
    .C(_13963_),
    .Y(_09509_));
 sky130_fd_sc_hd__a21oi_2 _23496_ (.A1(_13981_),
    .A2(_13971_),
    .B1(_13980_),
    .Y(_09510_));
 sky130_fd_sc_hd__o21ai_1 _23497_ (.A1(_09509_),
    .A2(_09508_),
    .B1(_09510_),
    .Y(_09511_));
 sky130_fd_sc_hd__nor3b_2 _23498_ (.A(_09493_),
    .B(_09508_),
    .C_N(_09488_),
    .Y(_09512_));
 sky130_fd_sc_hd__o21a_4 _23499_ (.A1(_09512_),
    .A2(_09511_),
    .B1(_13991_),
    .X(_09513_));
 sky130_fd_sc_hd__nor3_1 _23500_ (.A(_13991_),
    .B(_09511_),
    .C(_09512_),
    .Y(_09514_));
 sky130_fd_sc_hd__nor2_4 _23501_ (.A(_09513_),
    .B(_09514_),
    .Y(\hash.CA1.p3[15] ));
 sky130_fd_sc_hd__nor3_2 _23502_ (.A(_13954_),
    .B(_13963_),
    .C(_13990_),
    .Y(_09515_));
 sky130_fd_sc_hd__nand2_1 _23503_ (.A(_09510_),
    .B(_09515_),
    .Y(_09516_));
 sky130_fd_sc_hd__a21boi_2 _23504_ (.A1(_09510_),
    .A2(_09508_),
    .B1_N(_13991_),
    .Y(_09517_));
 sky130_fd_sc_hd__o22ai_1 _23505_ (.A1(_09501_),
    .A2(_09516_),
    .B1(_09517_),
    .B2(_13990_),
    .Y(_09518_));
 sky130_fd_sc_hd__xnor2_1 _23506_ (.A(_14000_),
    .B(_09518_),
    .Y(\hash.CA1.p3[16] ));
 sky130_fd_sc_hd__o21a_1 _23507_ (.A1(_14000_),
    .A2(_13999_),
    .B1(_14008_),
    .X(_09519_));
 sky130_fd_sc_hd__o31a_1 _23508_ (.A1(_13990_),
    .A2(_13999_),
    .A3(_09513_),
    .B1(_09519_),
    .X(_09520_));
 sky130_fd_sc_hd__o21ai_0 _23509_ (.A1(_13990_),
    .A2(_09513_),
    .B1(_14000_),
    .Y(_09521_));
 sky130_fd_sc_hd__nor3b_1 _23510_ (.A(_14008_),
    .B(_13999_),
    .C_N(_09521_),
    .Y(_09522_));
 sky130_fd_sc_hd__nor2_1 _23511_ (.A(_09520_),
    .B(_09522_),
    .Y(\hash.CA1.p3[17] ));
 sky130_fd_sc_hd__o221a_4 _23512_ (.A1(_09516_),
    .A2(_09501_),
    .B1(_09517_),
    .B2(_13990_),
    .C1(_14000_),
    .X(_09523_));
 sky130_fd_sc_hd__o21a_1 _23513_ (.A1(_13999_),
    .A2(_09523_),
    .B1(_14008_),
    .X(_09524_));
 sky130_fd_sc_hd__nor2_1 _23514_ (.A(_14007_),
    .B(_09524_),
    .Y(_09525_));
 sky130_fd_sc_hd__xnor2_1 _23515_ (.A(_14016_),
    .B(_09525_),
    .Y(\hash.CA1.p3[18] ));
 sky130_fd_sc_hd__o21a_1 _23516_ (.A1(_14007_),
    .A2(_09520_),
    .B1(_14016_),
    .X(_09526_));
 sky130_fd_sc_hd__nor2_1 _23517_ (.A(_14015_),
    .B(_09526_),
    .Y(_09527_));
 sky130_fd_sc_hd__xnor2_1 _23518_ (.A(_14024_),
    .B(_09527_),
    .Y(\hash.CA1.p3[19] ));
 sky130_fd_sc_hd__o21a_1 _23519_ (.A1(_14008_),
    .A2(_14007_),
    .B1(_14016_),
    .X(_09528_));
 sky130_fd_sc_hd__o31ai_4 _23520_ (.A1(_13999_),
    .A2(_09523_),
    .A3(_14007_),
    .B1(_09528_),
    .Y(_09529_));
 sky130_fd_sc_hd__nand2b_1 _23521_ (.A_N(_14015_),
    .B(_09529_),
    .Y(_09530_));
 sky130_fd_sc_hd__a21oi_1 _23522_ (.A1(_14024_),
    .A2(_09530_),
    .B1(_14023_),
    .Y(_09531_));
 sky130_fd_sc_hd__xnor2_1 _23523_ (.A(_14032_),
    .B(_09531_),
    .Y(\hash.CA1.p3[20] ));
 sky130_fd_sc_hd__or3_4 _23524_ (.A(_14007_),
    .B(_14015_),
    .C(_14023_),
    .X(_09532_));
 sky130_fd_sc_hd__or2_0 _23525_ (.A(_09532_),
    .B(_09520_),
    .X(_09533_));
 sky130_fd_sc_hd__or3_4 _23526_ (.A(_14016_),
    .B(_14015_),
    .C(_14023_),
    .X(_09534_));
 sky130_fd_sc_hd__or2_4 _23527_ (.A(_14024_),
    .B(_14023_),
    .X(_09535_));
 sky130_fd_sc_hd__a41o_1 _23528_ (.A1(_09533_),
    .A2(_14032_),
    .A3(_09534_),
    .A4(_09535_),
    .B1(_14031_),
    .X(_09536_));
 sky130_fd_sc_hd__xor2_1 _23529_ (.A(_14041_),
    .B(_09536_),
    .X(\hash.CA1.p3[21] ));
 sky130_fd_sc_hd__nor3_1 _23530_ (.A(_14015_),
    .B(_14023_),
    .C(_14031_),
    .Y(_09537_));
 sky130_fd_sc_hd__a21oi_1 _23531_ (.A1(_14032_),
    .A2(_09535_),
    .B1(_14031_),
    .Y(_09538_));
 sky130_fd_sc_hd__a21oi_2 _23532_ (.A1(_09537_),
    .A2(_09529_),
    .B1(_09538_),
    .Y(_09539_));
 sky130_fd_sc_hd__a21oi_1 _23533_ (.A1(_14041_),
    .A2(_09539_),
    .B1(_14040_),
    .Y(_09540_));
 sky130_fd_sc_hd__xnor2_1 _23534_ (.A(_14051_),
    .B(_09540_),
    .Y(\hash.CA1.p3[22] ));
 sky130_fd_sc_hd__and3_1 _23535_ (.A(_14032_),
    .B(_14041_),
    .C(_14051_),
    .X(_09541_));
 sky130_fd_sc_hd__o2111ai_2 _23536_ (.A1(_09520_),
    .A2(_09532_),
    .B1(_09534_),
    .C1(_09535_),
    .D1(_09541_),
    .Y(_09542_));
 sky130_fd_sc_hd__and3_1 _23537_ (.A(_14041_),
    .B(_14051_),
    .C(_14031_),
    .X(_09543_));
 sky130_fd_sc_hd__a21oi_1 _23538_ (.A1(_14051_),
    .A2(_14040_),
    .B1(_09543_),
    .Y(_09544_));
 sky130_fd_sc_hd__nand3b_1 _23539_ (.A_N(_14050_),
    .B(_09544_),
    .C(_09542_),
    .Y(_09545_));
 sky130_fd_sc_hd__xor2_1 _23540_ (.A(_14061_),
    .B(_09545_),
    .X(\hash.CA1.p3[23] ));
 sky130_fd_sc_hd__nand2_1 _23541_ (.A(_14061_),
    .B(_14050_),
    .Y(_09546_));
 sky130_fd_sc_hd__nand3_1 _23542_ (.A(_14051_),
    .B(_14061_),
    .C(_14040_),
    .Y(_09547_));
 sky130_fd_sc_hd__nand2_1 _23543_ (.A(_09546_),
    .B(_09547_),
    .Y(_09548_));
 sky130_fd_sc_hd__a41oi_2 _23544_ (.A1(_14041_),
    .A2(_14051_),
    .A3(_09539_),
    .A4(_14061_),
    .B1(_09548_),
    .Y(_09549_));
 sky130_fd_sc_hd__nor2b_4 _23545_ (.A(_14060_),
    .B_N(_09549_),
    .Y(_09550_));
 sky130_fd_sc_hd__xnor2_1 _23546_ (.A(_09550_),
    .B(_14071_),
    .Y(\hash.CA1.p3[24] ));
 sky130_fd_sc_hd__nor3_1 _23547_ (.A(_14050_),
    .B(_14060_),
    .C(_14070_),
    .Y(_09551_));
 sky130_fd_sc_hd__or2_0 _23548_ (.A(_14071_),
    .B(_14070_),
    .X(_09552_));
 sky130_fd_sc_hd__o31ai_1 _23549_ (.A1(_14061_),
    .A2(_14060_),
    .A3(_14070_),
    .B1(_09552_),
    .Y(_09553_));
 sky130_fd_sc_hd__a31o_4 _23550_ (.A1(_09544_),
    .A2(_09542_),
    .A3(_09551_),
    .B1(_09553_),
    .X(_09554_));
 sky130_fd_sc_hd__xnor2_2 _23551_ (.A(_14081_),
    .B(_09554_),
    .Y(\hash.CA1.p3[25] ));
 sky130_fd_sc_hd__nor3_2 _23552_ (.A(_14060_),
    .B(_14070_),
    .C(_14080_),
    .Y(_09555_));
 sky130_fd_sc_hd__a21oi_1 _23553_ (.A1(_14081_),
    .A2(_09552_),
    .B1(_14080_),
    .Y(_09556_));
 sky130_fd_sc_hd__a21oi_4 _23554_ (.A1(_09555_),
    .A2(_09549_),
    .B1(_09556_),
    .Y(_09557_));
 sky130_fd_sc_hd__xor2_1 _23555_ (.A(_14090_),
    .B(_09557_),
    .X(\hash.CA1.p3[26] ));
 sky130_fd_sc_hd__nand2_1 _23556_ (.A(_14081_),
    .B(_14090_),
    .Y(_09558_));
 sky130_fd_sc_hd__a21oi_1 _23557_ (.A1(_14090_),
    .A2(_14080_),
    .B1(_14089_),
    .Y(_09559_));
 sky130_fd_sc_hd__o21ai_4 _23558_ (.A1(_09554_),
    .A2(_09558_),
    .B1(_09559_),
    .Y(_09560_));
 sky130_fd_sc_hd__xor2_1 _23559_ (.A(_09560_),
    .B(_14099_),
    .X(\hash.CA1.p3[27] ));
 sky130_fd_sc_hd__a21o_1 _23560_ (.A1(_09557_),
    .A2(_14090_),
    .B1(_14089_),
    .X(_09561_));
 sky130_fd_sc_hd__a21oi_2 _23561_ (.A1(_09561_),
    .A2(_14099_),
    .B1(_14098_),
    .Y(_09562_));
 sky130_fd_sc_hd__xnor2_1 _23562_ (.A(_09562_),
    .B(_14109_),
    .Y(\hash.CA1.p3[28] ));
 sky130_fd_sc_hd__a21o_1 _23563_ (.A1(_09560_),
    .A2(_14099_),
    .B1(_14098_),
    .X(_09563_));
 sky130_fd_sc_hd__a21oi_2 _23564_ (.A1(_09563_),
    .A2(_14109_),
    .B1(_14108_),
    .Y(_09564_));
 sky130_fd_sc_hd__xnor2_1 _23565_ (.A(_09564_),
    .B(_14118_),
    .Y(\hash.CA1.p3[29] ));
 sky130_fd_sc_hd__nand2_2 _23566_ (.A(_09557_),
    .B(_14090_),
    .Y(_09565_));
 sky130_fd_sc_hd__nand3_1 _23567_ (.A(_14099_),
    .B(_14109_),
    .C(_14118_),
    .Y(_09566_));
 sky130_fd_sc_hd__a21o_1 _23568_ (.A1(_14099_),
    .A2(_14089_),
    .B1(_14098_),
    .X(_09567_));
 sky130_fd_sc_hd__a21o_1 _23569_ (.A1(_14109_),
    .A2(_09567_),
    .B1(_14108_),
    .X(_09568_));
 sky130_fd_sc_hd__a21oi_1 _23570_ (.A1(_14118_),
    .A2(_09568_),
    .B1(_14117_),
    .Y(_09569_));
 sky130_fd_sc_hd__o21ai_2 _23571_ (.A1(_09566_),
    .A2(_09565_),
    .B1(_09569_),
    .Y(_09570_));
 sky130_fd_sc_hd__xor2_1 _23572_ (.A(_09570_),
    .B(_14127_),
    .X(\hash.CA1.p3[30] ));
 sky130_fd_sc_hd__nor3b_1 _23573_ (.A(_09566_),
    .B(_12651_),
    .C_N(_14127_),
    .Y(_09571_));
 sky130_fd_sc_hd__a21o_1 _23574_ (.A1(_14109_),
    .A2(_14098_),
    .B1(_14108_),
    .X(_09572_));
 sky130_fd_sc_hd__a21o_1 _23575_ (.A1(_14118_),
    .A2(_09572_),
    .B1(_14117_),
    .X(_09573_));
 sky130_fd_sc_hd__nor4b_2 _23576_ (.A(_14126_),
    .B(_09573_),
    .C(_09560_),
    .D_N(_12651_),
    .Y(_09574_));
 sky130_fd_sc_hd__a21oi_1 _23577_ (.A1(_14127_),
    .A2(_09573_),
    .B1(_14126_),
    .Y(_09575_));
 sky130_fd_sc_hd__nand2b_1 _23578_ (.A_N(_09573_),
    .B(_09566_),
    .Y(_09576_));
 sky130_fd_sc_hd__a21oi_1 _23579_ (.A1(_14127_),
    .A2(_09576_),
    .B1(_14126_),
    .Y(_09577_));
 sky130_fd_sc_hd__nand2_1 _23580_ (.A(_12651_),
    .B(_09577_),
    .Y(_09578_));
 sky130_fd_sc_hd__o21ai_0 _23581_ (.A1(_12651_),
    .A2(_09575_),
    .B1(_09578_),
    .Y(_09579_));
 sky130_fd_sc_hd__a211o_1 _23582_ (.A1(_09560_),
    .A2(_09571_),
    .B1(_09579_),
    .C1(_09574_),
    .X(_09580_));
 sky130_fd_sc_hd__xnor2_1 _23583_ (.A(_09449_),
    .B(_09580_),
    .Y(\hash.CA1.p3[31] ));
 sky130_fd_sc_hd__xnor2_4 _23584_ (.A(_12892_),
    .B(_13883_),
    .Y(\hash.CA1.p3[3] ));
 sky130_fd_sc_hd__xnor2_4 _23585_ (.A(_13893_),
    .B(_09473_),
    .Y(\hash.CA1.p3[4] ));
 sky130_fd_sc_hd__nand2_1 _23586_ (.A(_09474_),
    .B(_09483_),
    .Y(_09581_));
 sky130_fd_sc_hd__nor2_1 _23587_ (.A(_13902_),
    .B(_09581_),
    .Y(_09582_));
 sky130_fd_sc_hd__nor2_4 _23588_ (.A(_09484_),
    .B(_09582_),
    .Y(\hash.CA1.p3[5] ));
 sky130_fd_sc_hd__xor2_4 _23589_ (.A(_13910_),
    .B(_09476_),
    .X(\hash.CA1.p3[6] ));
 sky130_fd_sc_hd__inv_1 _23590_ (.A(_09485_),
    .Y(_09583_));
 sky130_fd_sc_hd__a21oi_2 _23591_ (.A1(_13910_),
    .A2(_09583_),
    .B1(_13909_),
    .Y(_09584_));
 sky130_fd_sc_hd__xnor2_4 _23592_ (.A(_13918_),
    .B(_09584_),
    .Y(\hash.CA1.p3[7] ));
 sky130_fd_sc_hd__nor2_2 _23593_ (.A(_13917_),
    .B(_09478_),
    .Y(_09585_));
 sky130_fd_sc_hd__xnor2_4 _23594_ (.A(_13927_),
    .B(_09585_),
    .Y(\hash.CA1.p3[8] ));
 sky130_fd_sc_hd__nor3_1 _23595_ (.A(_13936_),
    .B(_13926_),
    .C(_09489_),
    .Y(_09586_));
 sky130_fd_sc_hd__nor2_4 _23596_ (.A(_09490_),
    .B(_09586_),
    .Y(\hash.CA1.p3[9] ));
 sky130_fd_sc_hd__xor2_1 _23597_ (.A(\hash.CA1.k_i2[31] ),
    .B(_12495_),
    .X(_09587_));
 sky130_fd_sc_hd__xnor2_1 _23598_ (.A(_06418_),
    .B(_09587_),
    .Y(_09588_));
 sky130_fd_sc_hd__xnor2_1 _23599_ (.A(\hash.CA1.w_i2[31] ),
    .B(_09588_),
    .Y(_09589_));
 sky130_fd_sc_hd__o21bai_1 _23600_ (.A1(_08034_),
    .A2(_08038_),
    .B1_N(_13825_),
    .Y(_09590_));
 sky130_fd_sc_hd__a21o_1 _23601_ (.A1(_13833_),
    .A2(_09590_),
    .B1(_13832_),
    .X(_09591_));
 sky130_fd_sc_hd__a21oi_1 _23602_ (.A1(_13839_),
    .A2(_09591_),
    .B1(_13838_),
    .Y(_09592_));
 sky130_fd_sc_hd__o21ai_0 _23603_ (.A1(_08035_),
    .A2(_08051_),
    .B1(_09592_),
    .Y(_09593_));
 sky130_fd_sc_hd__a21oi_1 _23604_ (.A1(_13844_),
    .A2(_09593_),
    .B1(_13843_),
    .Y(_09594_));
 sky130_fd_sc_hd__xnor2_1 _23605_ (.A(_09589_),
    .B(_09594_),
    .Y(\hash.CA1.p4[31] ));
 sky130_fd_sc_hd__inv_2 _23606_ (.A(_13723_),
    .Y(_09595_));
 sky130_fd_sc_hd__a21o_1 _23607_ (.A1(_13712_),
    .A2(_13704_),
    .B1(_13711_),
    .X(_09596_));
 sky130_fd_sc_hd__a21oi_2 _23608_ (.A1(_13718_),
    .A2(_09596_),
    .B1(_13717_),
    .Y(_09597_));
 sky130_fd_sc_hd__inv_1 _23609_ (.A(_13698_),
    .Y(_09598_));
 sky130_fd_sc_hd__clkinv_1 _23610_ (.A(_13680_),
    .Y(_09599_));
 sky130_fd_sc_hd__nor2b_1 _23611_ (.A(_12896_),
    .B_N(_13675_),
    .Y(_09600_));
 sky130_fd_sc_hd__o21ai_1 _23612_ (.A1(_13674_),
    .A2(_09600_),
    .B1(_13681_),
    .Y(_09601_));
 sky130_fd_sc_hd__a21boi_2 _23613_ (.A1(_09599_),
    .A2(_09601_),
    .B1_N(_13687_),
    .Y(_09602_));
 sky130_fd_sc_hd__o21a_4 _23614_ (.A1(_13686_),
    .A2(_09602_),
    .B1(_13693_),
    .X(_09603_));
 sky130_fd_sc_hd__o21ai_2 _23615_ (.A1(_13692_),
    .A2(_09603_),
    .B1(_13699_),
    .Y(_09604_));
 sky130_fd_sc_hd__and3_4 _23616_ (.A(_13705_),
    .B(_13712_),
    .C(_13718_),
    .X(_09605_));
 sky130_fd_sc_hd__a21bo_4 _23617_ (.A1(_09598_),
    .A2(_09604_),
    .B1_N(_09605_),
    .X(_09606_));
 sky130_fd_sc_hd__nand2_1 _23618_ (.A(_09597_),
    .B(_09606_),
    .Y(_09607_));
 sky130_fd_sc_hd__xnor2_1 _23619_ (.A(_09595_),
    .B(_09607_),
    .Y(\hash.CA1.p5[10] ));
 sky130_fd_sc_hd__inv_1 _23620_ (.A(_13681_),
    .Y(_09608_));
 sky130_fd_sc_hd__a21o_1 _23621_ (.A1(_12898_),
    .A2(_13670_),
    .B1(_13669_),
    .X(_09609_));
 sky130_fd_sc_hd__a21oi_2 _23622_ (.A1(_13675_),
    .A2(_09609_),
    .B1(_13674_),
    .Y(_09610_));
 sky130_fd_sc_hd__o21ai_2 _23623_ (.A1(_09608_),
    .A2(_09610_),
    .B1(_09599_),
    .Y(_09611_));
 sky130_fd_sc_hd__a21oi_4 _23624_ (.A1(_13687_),
    .A2(_09611_),
    .B1(_13686_),
    .Y(_09612_));
 sky130_fd_sc_hd__nor2_2 _23625_ (.A(_13692_),
    .B(_13698_),
    .Y(_09613_));
 sky130_fd_sc_hd__nand3_2 _23626_ (.A(_13723_),
    .B(_13729_),
    .C(_09605_),
    .Y(_09614_));
 sky130_fd_sc_hd__o21a_1 _23627_ (.A1(_13693_),
    .A2(_13692_),
    .B1(_13699_),
    .X(_09615_));
 sky130_fd_sc_hd__nor2_2 _23628_ (.A(_13698_),
    .B(_09615_),
    .Y(_09616_));
 sky130_fd_sc_hd__a211oi_4 _23629_ (.A1(_09612_),
    .A2(_09613_),
    .B1(_09614_),
    .C1(_09616_),
    .Y(_09617_));
 sky130_fd_sc_hd__nand2_1 _23630_ (.A(_13723_),
    .B(_13729_),
    .Y(_09618_));
 sky130_fd_sc_hd__nand2_1 _23631_ (.A(_13729_),
    .B(_13722_),
    .Y(_09619_));
 sky130_fd_sc_hd__o21ai_2 _23632_ (.A1(_09597_),
    .A2(_09618_),
    .B1(_09619_),
    .Y(_09620_));
 sky130_fd_sc_hd__a21oi_2 _23633_ (.A1(_09612_),
    .A2(_09613_),
    .B1(_09616_),
    .Y(_09621_));
 sky130_fd_sc_hd__nand2_1 _23634_ (.A(_09605_),
    .B(_09621_),
    .Y(_09622_));
 sky130_fd_sc_hd__nand2_1 _23635_ (.A(_09597_),
    .B(_09622_),
    .Y(_09623_));
 sky130_fd_sc_hd__a211oi_1 _23636_ (.A1(_13723_),
    .A2(_09623_),
    .B1(_13722_),
    .C1(_13729_),
    .Y(_09624_));
 sky130_fd_sc_hd__nor3_2 _23637_ (.A(_09617_),
    .B(_09620_),
    .C(_09624_),
    .Y(\hash.CA1.p5[11] ));
 sky130_fd_sc_hd__a21o_1 _23638_ (.A1(_13723_),
    .A2(_09607_),
    .B1(_13722_),
    .X(_09625_));
 sky130_fd_sc_hd__a21oi_2 _23639_ (.A1(_13729_),
    .A2(_09625_),
    .B1(_13728_),
    .Y(_09626_));
 sky130_fd_sc_hd__xnor2_2 _23640_ (.A(_13736_),
    .B(_09626_),
    .Y(\hash.CA1.p5[12] ));
 sky130_fd_sc_hd__o31ai_1 _23641_ (.A1(_13728_),
    .A2(_09617_),
    .A3(_09620_),
    .B1(_13736_),
    .Y(_09627_));
 sky130_fd_sc_hd__nand2b_2 _23642_ (.A_N(_13735_),
    .B(_09627_),
    .Y(_09628_));
 sky130_fd_sc_hd__xor2_2 _23643_ (.A(_13742_),
    .B(_09628_),
    .X(\hash.CA1.p5[13] ));
 sky130_fd_sc_hd__nand2_1 _23644_ (.A(_13729_),
    .B(_13736_),
    .Y(_09629_));
 sky130_fd_sc_hd__a211oi_2 _23645_ (.A1(_09597_),
    .A2(_09606_),
    .B1(_09629_),
    .C1(_09595_),
    .Y(_09630_));
 sky130_fd_sc_hd__nand2b_1 _23646_ (.A_N(_13728_),
    .B(_09619_),
    .Y(_09631_));
 sky130_fd_sc_hd__a21o_4 _23647_ (.A1(_13736_),
    .A2(_09631_),
    .B1(_13735_),
    .X(_09632_));
 sky130_fd_sc_hd__o21ai_1 _23648_ (.A1(_09630_),
    .A2(_09632_),
    .B1(_13742_),
    .Y(_09633_));
 sky130_fd_sc_hd__nand2b_4 _23649_ (.A_N(_13741_),
    .B(_09633_),
    .Y(_09634_));
 sky130_fd_sc_hd__xor2_1 _23650_ (.A(_13748_),
    .B(_09634_),
    .X(\hash.CA1.p5[14] ));
 sky130_fd_sc_hd__or3_1 _23651_ (.A(_13728_),
    .B(_13735_),
    .C(_13741_),
    .X(_09635_));
 sky130_fd_sc_hd__nor3_1 _23652_ (.A(_13736_),
    .B(_13735_),
    .C(_13741_),
    .Y(_09636_));
 sky130_fd_sc_hd__nor2_1 _23653_ (.A(_13742_),
    .B(_13741_),
    .Y(_09637_));
 sky130_fd_sc_hd__nor2_1 _23654_ (.A(_09636_),
    .B(_09637_),
    .Y(_09638_));
 sky130_fd_sc_hd__o31ai_2 _23655_ (.A1(_09617_),
    .A2(_09620_),
    .A3(_09635_),
    .B1(_09638_),
    .Y(_09639_));
 sky130_fd_sc_hd__nor2b_1 _23656_ (.A(_09639_),
    .B_N(_13748_),
    .Y(_09640_));
 sky130_fd_sc_hd__nor2_1 _23657_ (.A(_13747_),
    .B(_09640_),
    .Y(_09641_));
 sky130_fd_sc_hd__xnor2_1 _23658_ (.A(_13755_),
    .B(_09641_),
    .Y(\hash.CA1.p5[15] ));
 sky130_fd_sc_hd__a21o_1 _23659_ (.A1(_13748_),
    .A2(_09634_),
    .B1(_13747_),
    .X(_09642_));
 sky130_fd_sc_hd__a21o_4 _23660_ (.A1(_13755_),
    .A2(_09642_),
    .B1(_13754_),
    .X(_09643_));
 sky130_fd_sc_hd__xor2_1 _23661_ (.A(_13762_),
    .B(_09643_),
    .X(\hash.CA1.p5[16] ));
 sky130_fd_sc_hd__o21ai_0 _23662_ (.A1(_13747_),
    .A2(_09640_),
    .B1(_13755_),
    .Y(_09644_));
 sky130_fd_sc_hd__nand2b_1 _23663_ (.A_N(_13754_),
    .B(_09644_),
    .Y(_09645_));
 sky130_fd_sc_hd__a21oi_1 _23664_ (.A1(_13762_),
    .A2(_09645_),
    .B1(_13761_),
    .Y(_09646_));
 sky130_fd_sc_hd__xnor2_2 _23665_ (.A(_13769_),
    .B(_09646_),
    .Y(\hash.CA1.p5[17] ));
 sky130_fd_sc_hd__and2_4 _23666_ (.A(_13762_),
    .B(_13769_),
    .X(_09647_));
 sky130_fd_sc_hd__a221oi_1 _23667_ (.A1(_13769_),
    .A2(_13761_),
    .B1(_09643_),
    .B2(_09647_),
    .C1(_13768_),
    .Y(_09648_));
 sky130_fd_sc_hd__xnor2_1 _23668_ (.A(_13775_),
    .B(_09648_),
    .Y(\hash.CA1.p5[18] ));
 sky130_fd_sc_hd__clkinv_1 _23669_ (.A(_13780_),
    .Y(_09649_));
 sky130_fd_sc_hd__a21o_1 _23670_ (.A1(_13755_),
    .A2(_13747_),
    .B1(_13754_),
    .X(_09650_));
 sky130_fd_sc_hd__a21o_1 _23671_ (.A1(_13762_),
    .A2(_09650_),
    .B1(_13761_),
    .X(_09651_));
 sky130_fd_sc_hd__a21o_1 _23672_ (.A1(_13769_),
    .A2(_09651_),
    .B1(_13768_),
    .X(_09652_));
 sky130_fd_sc_hd__a21oi_1 _23673_ (.A1(_13775_),
    .A2(_09652_),
    .B1(_13774_),
    .Y(_09653_));
 sky130_fd_sc_hd__and4_4 _23674_ (.A(_13748_),
    .B(_13755_),
    .C(_13775_),
    .D(_09647_),
    .X(_09654_));
 sky130_fd_sc_hd__nand2b_1 _23675_ (.A_N(_09639_),
    .B(_09654_),
    .Y(_09655_));
 sky130_fd_sc_hd__nand2_1 _23676_ (.A(_09653_),
    .B(_09655_),
    .Y(_09656_));
 sky130_fd_sc_hd__xnor2_1 _23677_ (.A(_09649_),
    .B(_09656_),
    .Y(\hash.CA1.p5[19] ));
 sky130_fd_sc_hd__o21bai_1 _23678_ (.A1(_09649_),
    .A2(_09653_),
    .B1_N(_13779_),
    .Y(_09657_));
 sky130_fd_sc_hd__a31oi_1 _23679_ (.A1(_13780_),
    .A2(_09634_),
    .A3(_09654_),
    .B1(_09657_),
    .Y(_09658_));
 sky130_fd_sc_hd__xnor2_1 _23680_ (.A(_13785_),
    .B(_09658_),
    .Y(\hash.CA1.p5[20] ));
 sky130_fd_sc_hd__nand3_1 _23681_ (.A(_13780_),
    .B(_13785_),
    .C(_09654_),
    .Y(_09659_));
 sky130_fd_sc_hd__a21oi_1 _23682_ (.A1(_13785_),
    .A2(_09657_),
    .B1(_13784_),
    .Y(_09660_));
 sky130_fd_sc_hd__o21ai_2 _23683_ (.A1(_09639_),
    .A2(_09659_),
    .B1(_09660_),
    .Y(_09661_));
 sky130_fd_sc_hd__xor2_1 _23684_ (.A(_13790_),
    .B(_09661_),
    .X(\hash.CA1.p5[21] ));
 sky130_fd_sc_hd__o2111ai_2 _23685_ (.A1(_09630_),
    .A2(_09632_),
    .B1(_09654_),
    .C1(_13780_),
    .D1(_13742_),
    .Y(_09662_));
 sky130_fd_sc_hd__nor2_1 _23686_ (.A(_09649_),
    .B(_09653_),
    .Y(_09663_));
 sky130_fd_sc_hd__a31oi_2 _23687_ (.A1(_13780_),
    .A2(_13741_),
    .A3(_09654_),
    .B1(_09663_),
    .Y(_09664_));
 sky130_fd_sc_hd__nor3_1 _23688_ (.A(_13779_),
    .B(_13784_),
    .C(_13789_),
    .Y(_09665_));
 sky130_fd_sc_hd__or2_0 _23689_ (.A(_13785_),
    .B(_13784_),
    .X(_09666_));
 sky130_fd_sc_hd__a21oi_2 _23690_ (.A1(_13790_),
    .A2(_09666_),
    .B1(_13789_),
    .Y(_09667_));
 sky130_fd_sc_hd__a31oi_4 _23691_ (.A1(_09662_),
    .A2(_09664_),
    .A3(_09665_),
    .B1(_09667_),
    .Y(_09668_));
 sky130_fd_sc_hd__xor2_1 _23692_ (.A(_13795_),
    .B(_09668_),
    .X(\hash.CA1.p5[22] ));
 sky130_fd_sc_hd__inv_1 _23693_ (.A(_13801_),
    .Y(_09669_));
 sky130_fd_sc_hd__a21oi_1 _23694_ (.A1(_13795_),
    .A2(_13789_),
    .B1(_13794_),
    .Y(_09670_));
 sky130_fd_sc_hd__nand3_1 _23695_ (.A(_13790_),
    .B(_13795_),
    .C(_09661_),
    .Y(_09671_));
 sky130_fd_sc_hd__nand2_1 _23696_ (.A(_09670_),
    .B(_09671_),
    .Y(_09672_));
 sky130_fd_sc_hd__xnor2_1 _23697_ (.A(_09669_),
    .B(_09672_),
    .Y(\hash.CA1.p5[23] ));
 sky130_fd_sc_hd__a21o_1 _23698_ (.A1(_13795_),
    .A2(_09668_),
    .B1(_13794_),
    .X(_09673_));
 sky130_fd_sc_hd__a21oi_1 _23699_ (.A1(_13801_),
    .A2(_09673_),
    .B1(_13800_),
    .Y(_09674_));
 sky130_fd_sc_hd__xnor2_1 _23700_ (.A(_13808_),
    .B(_09674_),
    .Y(\hash.CA1.p5[24] ));
 sky130_fd_sc_hd__nand2_1 _23701_ (.A(_13801_),
    .B(_13808_),
    .Y(_09675_));
 sky130_fd_sc_hd__o21bai_1 _23702_ (.A1(_09669_),
    .A2(_09670_),
    .B1_N(_13800_),
    .Y(_09676_));
 sky130_fd_sc_hd__a21oi_1 _23703_ (.A1(_13808_),
    .A2(_09676_),
    .B1(_13807_),
    .Y(_09677_));
 sky130_fd_sc_hd__o21ai_0 _23704_ (.A1(_09671_),
    .A2(_09675_),
    .B1(_09677_),
    .Y(_09678_));
 sky130_fd_sc_hd__xor2_1 _23705_ (.A(_13815_),
    .B(_09678_),
    .X(\hash.CA1.p5[25] ));
 sky130_fd_sc_hd__and2_4 _23706_ (.A(_13801_),
    .B(_13808_),
    .X(_09679_));
 sky130_fd_sc_hd__nand4_1 _23707_ (.A(_13795_),
    .B(_13815_),
    .C(_09668_),
    .D(_09679_),
    .Y(_09680_));
 sky130_fd_sc_hd__a21oi_1 _23708_ (.A1(_13808_),
    .A2(_13800_),
    .B1(_13807_),
    .Y(_09681_));
 sky130_fd_sc_hd__nor2b_1 _23709_ (.A(_09681_),
    .B_N(_13815_),
    .Y(_09682_));
 sky130_fd_sc_hd__a31oi_1 _23710_ (.A1(_13815_),
    .A2(_13794_),
    .A3(_09679_),
    .B1(_09682_),
    .Y(_09683_));
 sky130_fd_sc_hd__nand2_1 _23711_ (.A(_09680_),
    .B(_09683_),
    .Y(_09684_));
 sky130_fd_sc_hd__nor2_1 _23712_ (.A(_13814_),
    .B(_09684_),
    .Y(_09685_));
 sky130_fd_sc_hd__xnor2_1 _23713_ (.A(_13822_),
    .B(_09685_),
    .Y(\hash.CA1.p5[26] ));
 sky130_fd_sc_hd__nand2_1 _23714_ (.A(_13790_),
    .B(_13795_),
    .Y(_09686_));
 sky130_fd_sc_hd__nand2_1 _23715_ (.A(_13815_),
    .B(_09679_),
    .Y(_09687_));
 sky130_fd_sc_hd__nor3b_1 _23716_ (.A(_09686_),
    .B(_09687_),
    .C_N(_09661_),
    .Y(_09688_));
 sky130_fd_sc_hd__nor2b_1 _23717_ (.A(_09677_),
    .B_N(_13815_),
    .Y(_09689_));
 sky130_fd_sc_hd__o31ai_1 _23718_ (.A1(_13814_),
    .A2(_09688_),
    .A3(_09689_),
    .B1(_13822_),
    .Y(_09690_));
 sky130_fd_sc_hd__nor2b_1 _23719_ (.A(_13821_),
    .B_N(_09690_),
    .Y(_09691_));
 sky130_fd_sc_hd__xnor2_1 _23720_ (.A(_13829_),
    .B(_09691_),
    .Y(\hash.CA1.p5[27] ));
 sky130_fd_sc_hd__nor3_1 _23721_ (.A(_13814_),
    .B(_13821_),
    .C(_13828_),
    .Y(_09692_));
 sky130_fd_sc_hd__or2_4 _23722_ (.A(_13829_),
    .B(_13828_),
    .X(_09693_));
 sky130_fd_sc_hd__o31ai_1 _23723_ (.A1(_13822_),
    .A2(_13821_),
    .A3(_13828_),
    .B1(_09693_),
    .Y(_09694_));
 sky130_fd_sc_hd__a31oi_1 _23724_ (.A1(_09680_),
    .A2(_09683_),
    .A3(_09692_),
    .B1(_09694_),
    .Y(_09695_));
 sky130_fd_sc_hd__xor2_1 _23725_ (.A(_13836_),
    .B(_09695_),
    .X(\hash.CA1.p5[28] ));
 sky130_fd_sc_hd__inv_1 _23726_ (.A(_13842_),
    .Y(_09696_));
 sky130_fd_sc_hd__nor3_1 _23727_ (.A(_13821_),
    .B(_13828_),
    .C(_13835_),
    .Y(_09697_));
 sky130_fd_sc_hd__a21oi_1 _23728_ (.A1(_13836_),
    .A2(_09693_),
    .B1(_13835_),
    .Y(_09698_));
 sky130_fd_sc_hd__a21oi_2 _23729_ (.A1(_09690_),
    .A2(_09697_),
    .B1(_09698_),
    .Y(_09699_));
 sky130_fd_sc_hd__xnor2_1 _23730_ (.A(_09696_),
    .B(_09699_),
    .Y(\hash.CA1.p5[29] ));
 sky130_fd_sc_hd__xnor2_1 _23731_ (.A(_12896_),
    .B(_13675_),
    .Y(\hash.CA1.p5[2] ));
 sky130_fd_sc_hd__a21oi_1 _23732_ (.A1(_13836_),
    .A2(_09695_),
    .B1(_13835_),
    .Y(_09700_));
 sky130_fd_sc_hd__o21bai_1 _23733_ (.A1(_09696_),
    .A2(_09700_),
    .B1_N(_13841_),
    .Y(_09701_));
 sky130_fd_sc_hd__xor2_1 _23734_ (.A(_13847_),
    .B(_09701_),
    .X(\hash.CA1.p5[30] ));
 sky130_fd_sc_hd__a21o_1 _23735_ (.A1(_13842_),
    .A2(_09699_),
    .B1(_13841_),
    .X(_09702_));
 sky130_fd_sc_hd__a21oi_1 _23736_ (.A1(_13847_),
    .A2(_09702_),
    .B1(_13846_),
    .Y(_09703_));
 sky130_fd_sc_hd__nand2_2 _23737_ (.A(_06002_),
    .B(\hash.CA2.a_dash[31] ),
    .Y(_09704_));
 sky130_fd_sc_hd__xnor2_1 _23738_ (.A(_09703_),
    .B(_09704_),
    .Y(_09705_));
 sky130_fd_sc_hd__xnor2_1 _23739_ (.A(\hash.CA1.p4[31] ),
    .B(_09705_),
    .Y(\hash.CA1.p5[31] ));
 sky130_fd_sc_hd__xnor2_1 _23740_ (.A(_13681_),
    .B(_09610_),
    .Y(\hash.CA1.p5[3] ));
 sky130_fd_sc_hd__nand2_1 _23741_ (.A(_09599_),
    .B(_09601_),
    .Y(_09706_));
 sky130_fd_sc_hd__nor2_1 _23742_ (.A(_13687_),
    .B(_09706_),
    .Y(_09707_));
 sky130_fd_sc_hd__nor2_1 _23743_ (.A(_09602_),
    .B(_09707_),
    .Y(\hash.CA1.p5[4] ));
 sky130_fd_sc_hd__xnor2_2 _23744_ (.A(_13693_),
    .B(_09612_),
    .Y(\hash.CA1.p5[5] ));
 sky130_fd_sc_hd__nor2_1 _23745_ (.A(_13692_),
    .B(_09603_),
    .Y(_09708_));
 sky130_fd_sc_hd__xnor2_2 _23746_ (.A(_13699_),
    .B(_09708_),
    .Y(\hash.CA1.p5[6] ));
 sky130_fd_sc_hd__xor2_1 _23747_ (.A(_13705_),
    .B(_09621_),
    .X(\hash.CA1.p5[7] ));
 sky130_fd_sc_hd__nand2_1 _23748_ (.A(_09598_),
    .B(_09604_),
    .Y(_09709_));
 sky130_fd_sc_hd__a21oi_1 _23749_ (.A1(_13705_),
    .A2(_09709_),
    .B1(_13704_),
    .Y(_09710_));
 sky130_fd_sc_hd__xnor2_1 _23750_ (.A(_13712_),
    .B(_09710_),
    .Y(\hash.CA1.p5[8] ));
 sky130_fd_sc_hd__inv_1 _23751_ (.A(_13712_),
    .Y(_09711_));
 sky130_fd_sc_hd__a21oi_1 _23752_ (.A1(_13705_),
    .A2(_09621_),
    .B1(_13704_),
    .Y(_09712_));
 sky130_fd_sc_hd__o21bai_1 _23753_ (.A1(_09711_),
    .A2(_09712_),
    .B1_N(_13711_),
    .Y(_09713_));
 sky130_fd_sc_hd__xor2_1 _23754_ (.A(_13718_),
    .B(_09713_),
    .X(\hash.CA1.p5[9] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_637 ();
 sky130_fd_sc_hd__or2_4 _23764_ (.A(\hash.CA2.b_dash[1] ),
    .B(net343),
    .X(_12657_));
 sky130_fd_sc_hd__inv_1 _23765_ (.A(_12657_),
    .Y(_00751_));
 sky130_fd_sc_hd__or2_4 _23766_ (.A(net340),
    .B(\hash.CA2.a_dash[1] ),
    .X(_12899_));
 sky130_fd_sc_hd__clkinv_1 _23767_ (.A(_12899_),
    .Y(_00721_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_636 ();
 sky130_fd_sc_hd__or2_4 _23769_ (.A(net340),
    .B(_12922_),
    .X(\hash.CA1.b[0] ));
 sky130_fd_sc_hd__inv_1 _23770_ (.A(\hash.CA1.b[0] ),
    .Y(_00690_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_634 ();
 sky130_fd_sc_hd__nand4_1 _23773_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(_13541_),
    .D(\count_2[5] ),
    .Y(_09726_));
 sky130_fd_sc_hd__or2_4 _23774_ (.A(\count_2[6] ),
    .B(_09726_),
    .X(_09727_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_633 ();
 sky130_fd_sc_hd__clkinv_2 _23776_ (.A(_09727_),
    .Y(_00128_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_631 ();
 sky130_fd_sc_hd__clkinv_16 _23779_ (.A(net780),
    .Y(_09731_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_627 ();
 sky130_fd_sc_hd__nor3_4 _23784_ (.A(\count_1[5] ),
    .B(\count_1[4] ),
    .C(\count_1[3] ),
    .Y(_09735_));
 sky130_fd_sc_hd__nand2_4 _23785_ (.A(_13528_),
    .B(_09735_),
    .Y(_09736_));
 sky130_fd_sc_hd__nand2_8 _23786_ (.A(_09731_),
    .B(_09736_),
    .Y(_00127_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_625 ();
 sky130_fd_sc_hd__nor3b_4 _23789_ (.A(\count_1[5] ),
    .B(\count_1[4] ),
    .C_N(\count_1[3] ),
    .Y(_09739_));
 sky130_fd_sc_hd__nand2_2 _23790_ (.A(_13531_),
    .B(_09739_),
    .Y(_09740_));
 sky130_fd_sc_hd__nand2_8 _23791_ (.A(_09731_),
    .B(_09740_),
    .Y(_00126_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_624 ();
 sky130_fd_sc_hd__nand2_2 _23793_ (.A(_13529_),
    .B(_09739_),
    .Y(_09742_));
 sky130_fd_sc_hd__nand2_8 _23794_ (.A(_09731_),
    .B(_09742_),
    .Y(_00125_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_623 ();
 sky130_fd_sc_hd__nand2_4 _23796_ (.A(_13533_),
    .B(_09739_),
    .Y(_09744_));
 sky130_fd_sc_hd__nand2_8 _23797_ (.A(_09731_),
    .B(_09744_),
    .Y(_00124_));
 sky130_fd_sc_hd__nor3b_4 _23798_ (.A(\count_1[5] ),
    .B(\count_1[3] ),
    .C_N(\count_1[4] ),
    .Y(_09745_));
 sky130_fd_sc_hd__nand2_2 _23799_ (.A(_13528_),
    .B(_09745_),
    .Y(_09746_));
 sky130_fd_sc_hd__nand2_8 _23800_ (.A(_09731_),
    .B(_09746_),
    .Y(_00123_));
 sky130_fd_sc_hd__nand2_2 _23801_ (.A(_13531_),
    .B(_09745_),
    .Y(_09747_));
 sky130_fd_sc_hd__nand2_8 _23802_ (.A(_09731_),
    .B(_09747_),
    .Y(_00122_));
 sky130_fd_sc_hd__nand2_2 _23803_ (.A(_13529_),
    .B(_09745_),
    .Y(_09748_));
 sky130_fd_sc_hd__nand2_8 _23804_ (.A(_09731_),
    .B(_09748_),
    .Y(_00121_));
 sky130_fd_sc_hd__nand2_2 _23805_ (.A(_13533_),
    .B(_09745_),
    .Y(_09749_));
 sky130_fd_sc_hd__nand2_8 _23806_ (.A(_09731_),
    .B(_09749_),
    .Y(_00120_));
 sky130_fd_sc_hd__nand2_1 _23807_ (.A(\count_1[4] ),
    .B(\count_1[3] ),
    .Y(_09750_));
 sky130_fd_sc_hd__nor2_4 _23808_ (.A(\count_1[5] ),
    .B(_09750_),
    .Y(_09751_));
 sky130_fd_sc_hd__nand2_2 _23809_ (.A(_13528_),
    .B(_09751_),
    .Y(_09752_));
 sky130_fd_sc_hd__nand2_8 _23810_ (.A(_09731_),
    .B(_09752_),
    .Y(_00119_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_621 ();
 sky130_fd_sc_hd__nand2_2 _23813_ (.A(_13531_),
    .B(_09751_),
    .Y(_09755_));
 sky130_fd_sc_hd__nand2_8 _23814_ (.A(_09731_),
    .B(_09755_),
    .Y(_00118_));
 sky130_fd_sc_hd__nand2_2 _23815_ (.A(_13529_),
    .B(_09751_),
    .Y(_09756_));
 sky130_fd_sc_hd__nand2_8 _23816_ (.A(_09731_),
    .B(_09756_),
    .Y(_00117_));
 sky130_fd_sc_hd__nand2_2 _23817_ (.A(_13531_),
    .B(_09735_),
    .Y(_09757_));
 sky130_fd_sc_hd__nand2_8 _23818_ (.A(_09731_),
    .B(_09757_),
    .Y(_00116_));
 sky130_fd_sc_hd__nand2_4 _23819_ (.A(_13533_),
    .B(_09751_),
    .Y(_09758_));
 sky130_fd_sc_hd__nand2_8 _23820_ (.A(_09731_),
    .B(_09758_),
    .Y(_00115_));
 sky130_fd_sc_hd__nor3b_4 _23821_ (.A(\count_1[4] ),
    .B(\count_1[3] ),
    .C_N(\count_1[5] ),
    .Y(_09759_));
 sky130_fd_sc_hd__nand2_4 _23822_ (.A(_13528_),
    .B(_09759_),
    .Y(_09760_));
 sky130_fd_sc_hd__nand2_8 _23823_ (.A(_09731_),
    .B(_09760_),
    .Y(_00114_));
 sky130_fd_sc_hd__nand2_2 _23824_ (.A(_13531_),
    .B(_09759_),
    .Y(_09761_));
 sky130_fd_sc_hd__nand2_8 _23825_ (.A(_09731_),
    .B(_09761_),
    .Y(_00113_));
 sky130_fd_sc_hd__nand2_4 _23826_ (.A(_13529_),
    .B(_09759_),
    .Y(_09762_));
 sky130_fd_sc_hd__nand2_8 _23827_ (.A(_09731_),
    .B(_09762_),
    .Y(_00112_));
 sky130_fd_sc_hd__nand2_4 _23828_ (.A(_13533_),
    .B(_09759_),
    .Y(_09763_));
 sky130_fd_sc_hd__nand2_8 _23829_ (.A(_09731_),
    .B(_09763_),
    .Y(_00111_));
 sky130_fd_sc_hd__and3b_4 _23830_ (.A_N(\count_1[4] ),
    .B(\count_1[3] ),
    .C(\count_1[5] ),
    .X(_09764_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_620 ();
 sky130_fd_sc_hd__nand2_4 _23832_ (.A(_13528_),
    .B(_09764_),
    .Y(_09766_));
 sky130_fd_sc_hd__nand2_8 _23833_ (.A(_09731_),
    .B(_09766_),
    .Y(_00110_));
 sky130_fd_sc_hd__nand2_4 _23834_ (.A(_13531_),
    .B(_09764_),
    .Y(_09767_));
 sky130_fd_sc_hd__nand2_8 _23835_ (.A(_09731_),
    .B(_09767_),
    .Y(_00109_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_619 ();
 sky130_fd_sc_hd__nand2_2 _23837_ (.A(_13529_),
    .B(_09764_),
    .Y(_09769_));
 sky130_fd_sc_hd__nand2_8 _23838_ (.A(_09731_),
    .B(_09769_),
    .Y(_00108_));
 sky130_fd_sc_hd__nand2_4 _23839_ (.A(_13533_),
    .B(_09764_),
    .Y(_09770_));
 sky130_fd_sc_hd__nand2_8 _23840_ (.A(_09731_),
    .B(_09770_),
    .Y(_00107_));
 sky130_fd_sc_hd__and3b_4 _23841_ (.A_N(\count_1[3] ),
    .B(\count_1[4] ),
    .C(\count_1[5] ),
    .X(_09771_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_618 ();
 sky130_fd_sc_hd__nand2_2 _23843_ (.A(_13528_),
    .B(_09771_),
    .Y(_09773_));
 sky130_fd_sc_hd__nand2_8 _23844_ (.A(_09731_),
    .B(_09773_),
    .Y(_00106_));
 sky130_fd_sc_hd__nand2_4 _23845_ (.A(_13529_),
    .B(_09735_),
    .Y(_09774_));
 sky130_fd_sc_hd__nand2_8 _23846_ (.A(_09731_),
    .B(_09774_),
    .Y(_00105_));
 sky130_fd_sc_hd__nand2_2 _23847_ (.A(_13531_),
    .B(_09771_),
    .Y(_09775_));
 sky130_fd_sc_hd__nand2_8 _23848_ (.A(_09731_),
    .B(_09775_),
    .Y(_00104_));
 sky130_fd_sc_hd__nand2_4 _23849_ (.A(_13529_),
    .B(_09771_),
    .Y(_09776_));
 sky130_fd_sc_hd__nand2_8 _23850_ (.A(_09731_),
    .B(_09776_),
    .Y(_00103_));
 sky130_fd_sc_hd__nand2_2 _23851_ (.A(_13533_),
    .B(_09771_),
    .Y(_09777_));
 sky130_fd_sc_hd__nand2_8 _23852_ (.A(_09731_),
    .B(_09777_),
    .Y(_00102_));
 sky130_fd_sc_hd__and3_4 _23853_ (.A(\count_1[5] ),
    .B(\count_1[4] ),
    .C(\count_1[3] ),
    .X(_09778_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_617 ();
 sky130_fd_sc_hd__nand2_2 _23855_ (.A(_13528_),
    .B(_09778_),
    .Y(_09780_));
 sky130_fd_sc_hd__nand2_8 _23856_ (.A(_09731_),
    .B(_09780_),
    .Y(_00101_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_614 ();
 sky130_fd_sc_hd__nor3b_4 _23860_ (.A(\count_2[4] ),
    .B(\count_2[5] ),
    .C_N(\count_2[3] ),
    .Y(_09784_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_613 ();
 sky130_fd_sc_hd__nand2_4 _23862_ (.A(_13539_),
    .B(net551),
    .Y(_09786_));
 sky130_fd_sc_hd__nand2_8 _23863_ (.A(_09731_),
    .B(_09786_),
    .Y(_00095_));
 sky130_fd_sc_hd__nand2_4 _23864_ (.A(_13531_),
    .B(_09778_),
    .Y(_09787_));
 sky130_fd_sc_hd__nand2_8 _23865_ (.A(_09731_),
    .B(_09787_),
    .Y(_00100_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_611 ();
 sky130_fd_sc_hd__nand2_2 _23868_ (.A(_13537_),
    .B(_09784_),
    .Y(_09790_));
 sky130_fd_sc_hd__nand2_8 _23869_ (.A(_09731_),
    .B(_09790_),
    .Y(_00094_));
 sky130_fd_sc_hd__nand2_4 _23870_ (.A(_13541_),
    .B(_09784_),
    .Y(_09791_));
 sky130_fd_sc_hd__nand2_8 _23871_ (.A(_09731_),
    .B(_09791_),
    .Y(_00093_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_610 ();
 sky130_fd_sc_hd__nand2b_4 _23873_ (.A_N(\count_2[3] ),
    .B(\count_2[4] ),
    .Y(_09793_));
 sky130_fd_sc_hd__nor2_4 _23874_ (.A(\count_2[5] ),
    .B(_09793_),
    .Y(_09794_));
 sky130_fd_sc_hd__nand2_4 _23875_ (.A(_13536_),
    .B(_09794_),
    .Y(_09795_));
 sky130_fd_sc_hd__nand2_8 _23876_ (.A(_09731_),
    .B(_09795_),
    .Y(_00092_));
 sky130_fd_sc_hd__nand2_2 _23877_ (.A(_13539_),
    .B(_09794_),
    .Y(_09796_));
 sky130_fd_sc_hd__nand2_8 _23878_ (.A(_09731_),
    .B(_09796_),
    .Y(_00091_));
 sky130_fd_sc_hd__nor3_4 _23879_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(\count_2[5] ),
    .Y(_09797_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_609 ();
 sky130_fd_sc_hd__nand2_2 _23881_ (.A(_13536_),
    .B(_09797_),
    .Y(_09799_));
 sky130_fd_sc_hd__nand2_8 _23882_ (.A(_09731_),
    .B(_09799_),
    .Y(_00090_));
 sky130_fd_sc_hd__nand2_2 _23883_ (.A(_13537_),
    .B(_09794_),
    .Y(_09800_));
 sky130_fd_sc_hd__nand2_8 _23884_ (.A(_09731_),
    .B(_09800_),
    .Y(_00089_));
 sky130_fd_sc_hd__nand2_2 _23885_ (.A(_13529_),
    .B(_09778_),
    .Y(_09801_));
 sky130_fd_sc_hd__nand2_8 _23886_ (.A(_09731_),
    .B(_09801_),
    .Y(_00099_));
 sky130_fd_sc_hd__inv_6 _23887_ (.A(\count_2[5] ),
    .Y(_09802_));
 sky130_fd_sc_hd__nand2_4 _23888_ (.A(_13541_),
    .B(_09802_),
    .Y(_09803_));
 sky130_fd_sc_hd__o21ai_4 _23889_ (.A1(_09793_),
    .A2(_09803_),
    .B1(_09731_),
    .Y(_00088_));
 sky130_fd_sc_hd__nand2_4 _23890_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .Y(_09804_));
 sky130_fd_sc_hd__nor2_4 _23891_ (.A(\count_2[5] ),
    .B(_09804_),
    .Y(_09805_));
 sky130_fd_sc_hd__nand2_2 _23892_ (.A(_13536_),
    .B(_09805_),
    .Y(_09806_));
 sky130_fd_sc_hd__nand2_8 _23893_ (.A(_09731_),
    .B(_09806_),
    .Y(_00087_));
 sky130_fd_sc_hd__nand2_4 _23894_ (.A(_13539_),
    .B(_09805_),
    .Y(_09807_));
 sky130_fd_sc_hd__nand2_8 _23895_ (.A(_09731_),
    .B(_09807_),
    .Y(_00086_));
 sky130_fd_sc_hd__nand2_2 _23896_ (.A(_13537_),
    .B(_09805_),
    .Y(_09808_));
 sky130_fd_sc_hd__nand2_8 _23897_ (.A(_09731_),
    .B(_09808_),
    .Y(_00085_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_608 ();
 sky130_fd_sc_hd__nand2_2 _23899_ (.A(_13541_),
    .B(_09805_),
    .Y(_09810_));
 sky130_fd_sc_hd__nand2_8 _23900_ (.A(_09731_),
    .B(_09810_),
    .Y(_00084_));
 sky130_fd_sc_hd__nor3_4 _23901_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(_09802_),
    .Y(_09811_));
 sky130_fd_sc_hd__nand2_2 _23902_ (.A(_13536_),
    .B(_09811_),
    .Y(_09812_));
 sky130_fd_sc_hd__nand2_8 _23903_ (.A(_09731_),
    .B(_09812_),
    .Y(_00083_));
 sky130_fd_sc_hd__nand2_4 _23904_ (.A(_13533_),
    .B(_09778_),
    .Y(_09813_));
 sky130_fd_sc_hd__nand2_8 _23905_ (.A(_09731_),
    .B(_09813_),
    .Y(_00098_));
 sky130_fd_sc_hd__nand2_4 _23906_ (.A(_13539_),
    .B(_09811_),
    .Y(_09814_));
 sky130_fd_sc_hd__nand2_8 _23907_ (.A(_09731_),
    .B(_09814_),
    .Y(_00082_));
 sky130_fd_sc_hd__nand2_4 _23908_ (.A(_13537_),
    .B(_09811_),
    .Y(_09815_));
 sky130_fd_sc_hd__nand2_8 _23909_ (.A(_09731_),
    .B(_09815_),
    .Y(_00081_));
 sky130_fd_sc_hd__nand2_4 _23910_ (.A(_13541_),
    .B(\count_2[5] ),
    .Y(_09816_));
 sky130_fd_sc_hd__o31ai_4 _23911_ (.A1(\count_2[4] ),
    .A2(\count_2[3] ),
    .A3(_09816_),
    .B1(_09731_),
    .Y(_00080_));
 sky130_fd_sc_hd__nand2_4 _23912_ (.A(_13539_),
    .B(_09797_),
    .Y(_09817_));
 sky130_fd_sc_hd__nand2_8 _23913_ (.A(_09731_),
    .B(_09817_),
    .Y(_00079_));
 sky130_fd_sc_hd__nor3b_4 _23914_ (.A(_09802_),
    .B(\count_2[4] ),
    .C_N(\count_2[3] ),
    .Y(_09818_));
 sky130_fd_sc_hd__nand2_4 _23915_ (.A(_13536_),
    .B(_09818_),
    .Y(_09819_));
 sky130_fd_sc_hd__nand2_8 _23916_ (.A(_09731_),
    .B(_09819_),
    .Y(_00078_));
 sky130_fd_sc_hd__nand2_4 _23917_ (.A(_13539_),
    .B(_09818_),
    .Y(_09820_));
 sky130_fd_sc_hd__nand2_8 _23918_ (.A(_09731_),
    .B(_09820_),
    .Y(_00077_));
 sky130_fd_sc_hd__nand2_4 _23919_ (.A(_13533_),
    .B(_09735_),
    .Y(_09821_));
 sky130_fd_sc_hd__nand2_8 _23920_ (.A(_09731_),
    .B(_09821_),
    .Y(_00097_));
 sky130_fd_sc_hd__nand2_2 _23921_ (.A(_13537_),
    .B(_09818_),
    .Y(_09822_));
 sky130_fd_sc_hd__nand2_8 _23922_ (.A(_09731_),
    .B(_09822_),
    .Y(_00076_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_607 ();
 sky130_fd_sc_hd__nand2_2 _23924_ (.A(_13541_),
    .B(_09818_),
    .Y(_09824_));
 sky130_fd_sc_hd__nand2_8 _23925_ (.A(_09731_),
    .B(_09824_),
    .Y(_00075_));
 sky130_fd_sc_hd__nor2_4 _23926_ (.A(_09802_),
    .B(_09793_),
    .Y(_09825_));
 sky130_fd_sc_hd__nand2_2 _23927_ (.A(_13536_),
    .B(_09825_),
    .Y(_09826_));
 sky130_fd_sc_hd__nand2_8 _23928_ (.A(_09731_),
    .B(_09826_),
    .Y(_00074_));
 sky130_fd_sc_hd__nand2_4 _23929_ (.A(_13539_),
    .B(_09825_),
    .Y(_09827_));
 sky130_fd_sc_hd__nand2_8 _23930_ (.A(_09731_),
    .B(_09827_),
    .Y(_00073_));
 sky130_fd_sc_hd__nand2_4 _23931_ (.A(_13537_),
    .B(_09825_),
    .Y(_09828_));
 sky130_fd_sc_hd__nand2_8 _23932_ (.A(_09731_),
    .B(_09828_),
    .Y(_00072_));
 sky130_fd_sc_hd__o21ai_4 _23933_ (.A1(_09816_),
    .A2(_09793_),
    .B1(_09731_),
    .Y(_00071_));
 sky130_fd_sc_hd__nand2_2 _23934_ (.A(_13528_),
    .B(_09739_),
    .Y(_09829_));
 sky130_fd_sc_hd__nand2_8 _23935_ (.A(_09731_),
    .B(_09829_),
    .Y(_00096_));
 sky130_fd_sc_hd__nor2_4 _23936_ (.A(_09802_),
    .B(_09804_),
    .Y(_09830_));
 sky130_fd_sc_hd__nand2_2 _23937_ (.A(_13536_),
    .B(_09830_),
    .Y(_09831_));
 sky130_fd_sc_hd__nand2_8 _23938_ (.A(_09731_),
    .B(_09831_),
    .Y(_00070_));
 sky130_fd_sc_hd__nand2_2 _23939_ (.A(_13539_),
    .B(_09830_),
    .Y(_09832_));
 sky130_fd_sc_hd__nand2_8 _23940_ (.A(_09731_),
    .B(_09832_),
    .Y(_00069_));
 sky130_fd_sc_hd__nand2_4 _23941_ (.A(_13537_),
    .B(_09797_),
    .Y(_09833_));
 sky130_fd_sc_hd__nand2_8 _23942_ (.A(_09731_),
    .B(_09833_),
    .Y(_00068_));
 sky130_fd_sc_hd__nand2_4 _23943_ (.A(_13537_),
    .B(_09830_),
    .Y(_09834_));
 sky130_fd_sc_hd__nand2_8 _23944_ (.A(_09731_),
    .B(_09834_),
    .Y(_00067_));
 sky130_fd_sc_hd__nand2_8 _23945_ (.A(_09731_),
    .B(_09726_),
    .Y(_00066_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_606 ();
 sky130_fd_sc_hd__nor3_4 _23947_ (.A(\count_2[4] ),
    .B(\count_2[3] ),
    .C(_09803_),
    .Y(_09836_));
 sky130_fd_sc_hd__or2_4 _23948_ (.A(net1039),
    .B(_09836_),
    .X(_00065_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_605 ();
 sky130_fd_sc_hd__nand2_4 _23950_ (.A(_13536_),
    .B(net551),
    .Y(_09838_));
 sky130_fd_sc_hd__nand2_8 _23951_ (.A(_09731_),
    .B(_09838_),
    .Y(_00064_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_600 ();
 sky130_fd_sc_hd__mux4_2 _23957_ (.A0(\w[19][0] ),
    .A1(\w[17][0] ),
    .A2(\w[23][0] ),
    .A3(\w[21][0] ),
    .S0(net359),
    .S1(net309),
    .X(_09844_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_598 ();
 sky130_fd_sc_hd__mux4_2 _23960_ (.A0(\w[27][0] ),
    .A1(\w[25][0] ),
    .A2(\w[31][0] ),
    .A3(\w[29][0] ),
    .S0(net359),
    .S1(net309),
    .X(_09847_));
 sky130_fd_sc_hd__mux4_2 _23961_ (.A0(\w[3][0] ),
    .A1(\w[1][0] ),
    .A2(\w[7][0] ),
    .A3(\w[5][0] ),
    .S0(net359),
    .S1(net309),
    .X(_09848_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_595 ();
 sky130_fd_sc_hd__mux4_2 _23965_ (.A0(\w[11][0] ),
    .A1(\w[9][0] ),
    .A2(\w[15][0] ),
    .A3(\w[13][0] ),
    .S0(net359),
    .S1(net309),
    .X(_09852_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_594 ();
 sky130_fd_sc_hd__xor2_4 _23967_ (.A(\count_hash2[3] ),
    .B(_12908_),
    .X(_09854_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_593 ();
 sky130_fd_sc_hd__nand3_4 _23969_ (.A(\count_hash2[3] ),
    .B(\count_hash2[2] ),
    .C(\count_hash2[1] ),
    .Y(_09856_));
 sky130_fd_sc_hd__xor2_4 _23970_ (.A(\count_hash2[4] ),
    .B(_09856_),
    .X(_09857_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_592 ();
 sky130_fd_sc_hd__mux4_2 _23972_ (.A0(_09844_),
    .A1(_09847_),
    .A2(_09848_),
    .A3(_09852_),
    .S0(net333),
    .S1(net327),
    .X(_09859_));
 sky130_fd_sc_hd__mux4_2 _23973_ (.A0(\w[51][0] ),
    .A1(\w[49][0] ),
    .A2(\w[55][0] ),
    .A3(\w[53][0] ),
    .S0(net358),
    .S1(net310),
    .X(_09860_));
 sky130_fd_sc_hd__mux4_2 _23974_ (.A0(\w[59][0] ),
    .A1(\w[57][0] ),
    .A2(\w[63][0] ),
    .A3(\w[61][0] ),
    .S0(net358),
    .S1(net310),
    .X(_09861_));
 sky130_fd_sc_hd__mux4_2 _23975_ (.A0(\w[35][0] ),
    .A1(\w[33][0] ),
    .A2(\w[39][0] ),
    .A3(\w[37][0] ),
    .S0(net358),
    .S1(net310),
    .X(_09862_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_591 ();
 sky130_fd_sc_hd__mux4_2 _23977_ (.A0(\w[43][0] ),
    .A1(\w[41][0] ),
    .A2(\w[47][0] ),
    .A3(\w[45][0] ),
    .S0(net358),
    .S1(net310),
    .X(_09864_));
 sky130_fd_sc_hd__mux4_2 _23978_ (.A0(_09860_),
    .A1(_09861_),
    .A2(_09862_),
    .A3(_09864_),
    .S0(net336),
    .S1(net326),
    .X(_09865_));
 sky130_fd_sc_hd__nand3_4 _23979_ (.A(\count_hash2[4] ),
    .B(\count_hash2[3] ),
    .C(_12908_),
    .Y(_09866_));
 sky130_fd_sc_hd__xnor2_4 _23980_ (.A(\count_hash2[5] ),
    .B(_09866_),
    .Y(_09867_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_589 ();
 sky130_fd_sc_hd__mux2i_1 _23983_ (.A0(_09859_),
    .A1(_09865_),
    .S(net292),
    .Y(_09870_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_587 ();
 sky130_fd_sc_hd__nand4_1 _23986_ (.A(\count_hash1[4] ),
    .B(\count_hash1[3] ),
    .C(\count_hash1[5] ),
    .D(\count_hash1[2] ),
    .Y(_09873_));
 sky130_fd_sc_hd__nor2_2 _23987_ (.A(_12914_),
    .B(_09873_),
    .Y(_09874_));
 sky130_fd_sc_hd__or3_4 _23988_ (.A(\count_hash1[6] ),
    .B(net349),
    .C(_09874_),
    .X(_09875_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_584 ();
 sky130_fd_sc_hd__nand2_2 _23992_ (.A(net347),
    .B(\w[1][0] ),
    .Y(_09879_));
 sky130_fd_sc_hd__o21ai_4 _23993_ (.A1(_09870_),
    .A2(net285),
    .B1(_09879_),
    .Y(_00032_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_580 ();
 sky130_fd_sc_hd__mux4_2 _23998_ (.A0(\w[19][1] ),
    .A1(\w[17][1] ),
    .A2(\w[23][1] ),
    .A3(\w[21][1] ),
    .S0(net358),
    .S1(net310),
    .X(_09884_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_578 ();
 sky130_fd_sc_hd__mux4_2 _24001_ (.A0(\w[27][1] ),
    .A1(\w[25][1] ),
    .A2(\w[31][1] ),
    .A3(\w[29][1] ),
    .S0(net358),
    .S1(net310),
    .X(_09887_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_576 ();
 sky130_fd_sc_hd__mux4_2 _24004_ (.A0(\w[3][1] ),
    .A1(\w[1][1] ),
    .A2(\w[7][1] ),
    .A3(\w[5][1] ),
    .S0(net358),
    .S1(net310),
    .X(_09890_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_574 ();
 sky130_fd_sc_hd__mux4_2 _24007_ (.A0(\w[11][1] ),
    .A1(\w[9][1] ),
    .A2(\w[15][1] ),
    .A3(\w[13][1] ),
    .S0(net358),
    .S1(net310),
    .X(_09893_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_572 ();
 sky130_fd_sc_hd__mux4_2 _24010_ (.A0(_09884_),
    .A1(_09887_),
    .A2(_09890_),
    .A3(_09893_),
    .S0(net336),
    .S1(net326),
    .X(_09896_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_570 ();
 sky130_fd_sc_hd__mux4_2 _24013_ (.A0(\w[51][1] ),
    .A1(\w[49][1] ),
    .A2(\w[55][1] ),
    .A3(\w[53][1] ),
    .S0(net358),
    .S1(net310),
    .X(_09899_));
 sky130_fd_sc_hd__mux4_2 _24014_ (.A0(\w[59][1] ),
    .A1(\w[57][1] ),
    .A2(\w[63][1] ),
    .A3(\w[61][1] ),
    .S0(net358),
    .S1(net310),
    .X(_09900_));
 sky130_fd_sc_hd__mux4_2 _24015_ (.A0(\w[35][1] ),
    .A1(\w[33][1] ),
    .A2(\w[39][1] ),
    .A3(\w[37][1] ),
    .S0(net358),
    .S1(net310),
    .X(_09901_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_568 ();
 sky130_fd_sc_hd__mux4_2 _24018_ (.A0(\w[43][1] ),
    .A1(\w[41][1] ),
    .A2(\w[47][1] ),
    .A3(\w[45][1] ),
    .S0(net358),
    .S1(net310),
    .X(_09904_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_565 ();
 sky130_fd_sc_hd__mux4_2 _24022_ (.A0(_09899_),
    .A1(_09900_),
    .A2(_09901_),
    .A3(_09904_),
    .S0(net336),
    .S1(net326),
    .X(_09908_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_564 ();
 sky130_fd_sc_hd__mux2i_1 _24024_ (.A0(_09896_),
    .A1(_09908_),
    .S(net292),
    .Y(_09910_));
 sky130_fd_sc_hd__nand2_2 _24025_ (.A(net347),
    .B(\w[1][1] ),
    .Y(_09911_));
 sky130_fd_sc_hd__o21ai_4 _24026_ (.A1(net285),
    .A2(_09910_),
    .B1(_09911_),
    .Y(_00043_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_563 ();
 sky130_fd_sc_hd__mux4_2 _24028_ (.A0(\w[19][2] ),
    .A1(\w[17][2] ),
    .A2(\w[23][2] ),
    .A3(\w[21][2] ),
    .S0(net359),
    .S1(net309),
    .X(_09913_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_562 ();
 sky130_fd_sc_hd__mux4_2 _24030_ (.A0(\w[27][2] ),
    .A1(\w[25][2] ),
    .A2(\w[31][2] ),
    .A3(\w[29][2] ),
    .S0(net359),
    .S1(net309),
    .X(_09915_));
 sky130_fd_sc_hd__mux4_2 _24031_ (.A0(\w[3][2] ),
    .A1(\w[1][2] ),
    .A2(\w[7][2] ),
    .A3(\w[5][2] ),
    .S0(net359),
    .S1(net309),
    .X(_09916_));
 sky130_fd_sc_hd__mux4_2 _24032_ (.A0(\w[11][2] ),
    .A1(\w[9][2] ),
    .A2(\w[15][2] ),
    .A3(\w[13][2] ),
    .S0(net359),
    .S1(net309),
    .X(_09917_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_561 ();
 sky130_fd_sc_hd__mux4_2 _24034_ (.A0(_09913_),
    .A1(_09915_),
    .A2(_09916_),
    .A3(_09917_),
    .S0(net334),
    .S1(net327),
    .X(_09919_));
 sky130_fd_sc_hd__mux4_2 _24035_ (.A0(\w[51][2] ),
    .A1(\w[49][2] ),
    .A2(\w[55][2] ),
    .A3(\w[53][2] ),
    .S0(net362),
    .S1(net309),
    .X(_09920_));
 sky130_fd_sc_hd__mux4_2 _24036_ (.A0(\w[59][2] ),
    .A1(\w[57][2] ),
    .A2(\w[63][2] ),
    .A3(\w[61][2] ),
    .S0(net362),
    .S1(net309),
    .X(_09921_));
 sky130_fd_sc_hd__mux4_2 _24037_ (.A0(\w[35][2] ),
    .A1(\w[33][2] ),
    .A2(\w[39][2] ),
    .A3(\w[37][2] ),
    .S0(net362),
    .S1(net309),
    .X(_09922_));
 sky130_fd_sc_hd__mux4_2 _24038_ (.A0(\w[43][2] ),
    .A1(\w[41][2] ),
    .A2(\w[47][2] ),
    .A3(\w[45][2] ),
    .S0(net362),
    .S1(net309),
    .X(_09923_));
 sky130_fd_sc_hd__mux4_2 _24039_ (.A0(_09920_),
    .A1(_09921_),
    .A2(_09922_),
    .A3(_09923_),
    .S0(net336),
    .S1(net326),
    .X(_09924_));
 sky130_fd_sc_hd__mux2i_1 _24040_ (.A0(_09919_),
    .A1(_09924_),
    .S(net292),
    .Y(_09925_));
 sky130_fd_sc_hd__nand2_2 _24041_ (.A(net347),
    .B(\w[1][2] ),
    .Y(_09926_));
 sky130_fd_sc_hd__o21ai_4 _24042_ (.A1(net285),
    .A2(_09925_),
    .B1(_09926_),
    .Y(_00054_));
 sky130_fd_sc_hd__mux4_2 _24043_ (.A0(\w[19][3] ),
    .A1(\w[17][3] ),
    .A2(\w[23][3] ),
    .A3(\w[21][3] ),
    .S0(net358),
    .S1(net310),
    .X(_09927_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_560 ();
 sky130_fd_sc_hd__mux4_2 _24045_ (.A0(\w[27][3] ),
    .A1(\w[25][3] ),
    .A2(\w[31][3] ),
    .A3(\w[29][3] ),
    .S0(net358),
    .S1(net310),
    .X(_09929_));
 sky130_fd_sc_hd__mux4_2 _24046_ (.A0(\w[3][3] ),
    .A1(\w[1][3] ),
    .A2(\w[7][3] ),
    .A3(\w[5][3] ),
    .S0(net358),
    .S1(net310),
    .X(_09930_));
 sky130_fd_sc_hd__mux4_2 _24047_ (.A0(\w[11][3] ),
    .A1(\w[9][3] ),
    .A2(\w[15][3] ),
    .A3(\w[13][3] ),
    .S0(net358),
    .S1(net310),
    .X(_09931_));
 sky130_fd_sc_hd__mux4_2 _24048_ (.A0(_09927_),
    .A1(_09929_),
    .A2(_09930_),
    .A3(_09931_),
    .S0(net336),
    .S1(net326),
    .X(_09932_));
 sky130_fd_sc_hd__mux4_2 _24049_ (.A0(\w[51][3] ),
    .A1(\w[49][3] ),
    .A2(\w[55][3] ),
    .A3(\w[53][3] ),
    .S0(net360),
    .S1(net308),
    .X(_09933_));
 sky130_fd_sc_hd__mux4_2 _24050_ (.A0(\w[59][3] ),
    .A1(\w[57][3] ),
    .A2(\w[63][3] ),
    .A3(\w[61][3] ),
    .S0(net360),
    .S1(net308),
    .X(_09934_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_559 ();
 sky130_fd_sc_hd__mux4_2 _24052_ (.A0(\w[35][3] ),
    .A1(\w[33][3] ),
    .A2(\w[39][3] ),
    .A3(\w[37][3] ),
    .S0(net360),
    .S1(net308),
    .X(_09936_));
 sky130_fd_sc_hd__mux4_2 _24053_ (.A0(\w[43][3] ),
    .A1(\w[41][3] ),
    .A2(\w[47][3] ),
    .A3(\w[45][3] ),
    .S0(net360),
    .S1(net308),
    .X(_09937_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_558 ();
 sky130_fd_sc_hd__mux4_2 _24055_ (.A0(_09933_),
    .A1(_09934_),
    .A2(_09936_),
    .A3(_09937_),
    .S0(net335),
    .S1(net330),
    .X(_09939_));
 sky130_fd_sc_hd__mux2i_1 _24056_ (.A0(_09932_),
    .A1(_09939_),
    .S(net292),
    .Y(_09940_));
 sky130_fd_sc_hd__nand2_2 _24057_ (.A(net347),
    .B(\w[1][3] ),
    .Y(_09941_));
 sky130_fd_sc_hd__o21ai_4 _24058_ (.A1(net285),
    .A2(_09940_),
    .B1(_09941_),
    .Y(_00057_));
 sky130_fd_sc_hd__mux4_2 _24059_ (.A0(\w[19][4] ),
    .A1(\w[17][4] ),
    .A2(\w[23][4] ),
    .A3(\w[21][4] ),
    .S0(net359),
    .S1(net309),
    .X(_09942_));
 sky130_fd_sc_hd__mux4_2 _24060_ (.A0(\w[27][4] ),
    .A1(\w[25][4] ),
    .A2(\w[31][4] ),
    .A3(\w[29][4] ),
    .S0(net359),
    .S1(net309),
    .X(_09943_));
 sky130_fd_sc_hd__mux4_2 _24061_ (.A0(\w[3][4] ),
    .A1(\w[1][4] ),
    .A2(\w[7][4] ),
    .A3(\w[5][4] ),
    .S0(net359),
    .S1(net309),
    .X(_09944_));
 sky130_fd_sc_hd__mux4_2 _24062_ (.A0(\w[11][4] ),
    .A1(\w[9][4] ),
    .A2(\w[15][4] ),
    .A3(\w[13][4] ),
    .S0(net359),
    .S1(net309),
    .X(_09945_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_557 ();
 sky130_fd_sc_hd__mux4_2 _24064_ (.A0(_09942_),
    .A1(_09943_),
    .A2(_09944_),
    .A3(_09945_),
    .S0(net333),
    .S1(net327),
    .X(_09947_));
 sky130_fd_sc_hd__mux4_2 _24065_ (.A0(\w[51][4] ),
    .A1(\w[49][4] ),
    .A2(\w[55][4] ),
    .A3(\w[53][4] ),
    .S0(net358),
    .S1(net310),
    .X(_09948_));
 sky130_fd_sc_hd__mux4_2 _24066_ (.A0(\w[59][4] ),
    .A1(\w[57][4] ),
    .A2(\w[63][4] ),
    .A3(\w[61][4] ),
    .S0(net362),
    .S1(net310),
    .X(_09949_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_556 ();
 sky130_fd_sc_hd__mux4_2 _24068_ (.A0(\w[35][4] ),
    .A1(\w[33][4] ),
    .A2(\w[39][4] ),
    .A3(\w[37][4] ),
    .S0(net362),
    .S1(net310),
    .X(_09951_));
 sky130_fd_sc_hd__mux4_2 _24069_ (.A0(\w[43][4] ),
    .A1(\w[41][4] ),
    .A2(\w[47][4] ),
    .A3(\w[45][4] ),
    .S0(net358),
    .S1(net310),
    .X(_09952_));
 sky130_fd_sc_hd__mux4_2 _24070_ (.A0(_09948_),
    .A1(_09949_),
    .A2(_09951_),
    .A3(_09952_),
    .S0(net335),
    .S1(net328),
    .X(_09953_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_553 ();
 sky130_fd_sc_hd__mux2i_1 _24074_ (.A0(_09947_),
    .A1(_09953_),
    .S(net292),
    .Y(_09957_));
 sky130_fd_sc_hd__nand2_2 _24075_ (.A(net347),
    .B(\w[1][4] ),
    .Y(_09958_));
 sky130_fd_sc_hd__o21ai_4 _24076_ (.A1(net285),
    .A2(_09957_),
    .B1(_09958_),
    .Y(_00058_));
 sky130_fd_sc_hd__mux4_2 _24077_ (.A0(\w[19][5] ),
    .A1(\w[17][5] ),
    .A2(\w[23][5] ),
    .A3(\w[21][5] ),
    .S0(net358),
    .S1(net310),
    .X(_09959_));
 sky130_fd_sc_hd__mux4_2 _24078_ (.A0(\w[27][5] ),
    .A1(\w[25][5] ),
    .A2(\w[31][5] ),
    .A3(\w[29][5] ),
    .S0(net358),
    .S1(net310),
    .X(_09960_));
 sky130_fd_sc_hd__mux4_2 _24079_ (.A0(\w[3][5] ),
    .A1(\w[1][5] ),
    .A2(\w[7][5] ),
    .A3(\w[5][5] ),
    .S0(net358),
    .S1(net310),
    .X(_09961_));
 sky130_fd_sc_hd__mux4_2 _24080_ (.A0(\w[11][5] ),
    .A1(\w[9][5] ),
    .A2(\w[15][5] ),
    .A3(\w[13][5] ),
    .S0(net358),
    .S1(net310),
    .X(_09962_));
 sky130_fd_sc_hd__mux4_2 _24081_ (.A0(_09959_),
    .A1(_09960_),
    .A2(_09961_),
    .A3(_09962_),
    .S0(net333),
    .S1(net326),
    .X(_09963_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_552 ();
 sky130_fd_sc_hd__mux4_2 _24083_ (.A0(\w[51][5] ),
    .A1(\w[49][5] ),
    .A2(\w[55][5] ),
    .A3(\w[53][5] ),
    .S0(net360),
    .S1(net308),
    .X(_09965_));
 sky130_fd_sc_hd__mux4_2 _24084_ (.A0(\w[59][5] ),
    .A1(\w[57][5] ),
    .A2(\w[63][5] ),
    .A3(\w[61][5] ),
    .S0(net360),
    .S1(net308),
    .X(_09966_));
 sky130_fd_sc_hd__mux4_2 _24085_ (.A0(\w[35][5] ),
    .A1(\w[33][5] ),
    .A2(\w[39][5] ),
    .A3(\w[37][5] ),
    .S0(net360),
    .S1(net308),
    .X(_09967_));
 sky130_fd_sc_hd__mux4_2 _24086_ (.A0(\w[43][5] ),
    .A1(\w[41][5] ),
    .A2(\w[47][5] ),
    .A3(\w[45][5] ),
    .S0(net360),
    .S1(net308),
    .X(_09968_));
 sky130_fd_sc_hd__mux4_2 _24087_ (.A0(_09965_),
    .A1(_09966_),
    .A2(_09967_),
    .A3(_09968_),
    .S0(net335),
    .S1(net330),
    .X(_09969_));
 sky130_fd_sc_hd__mux2i_1 _24088_ (.A0(_09963_),
    .A1(_09969_),
    .S(net292),
    .Y(_09970_));
 sky130_fd_sc_hd__nand2_2 _24089_ (.A(net347),
    .B(\w[1][5] ),
    .Y(_09971_));
 sky130_fd_sc_hd__o21ai_4 _24090_ (.A1(net285),
    .A2(_09970_),
    .B1(_09971_),
    .Y(_00059_));
 sky130_fd_sc_hd__mux4_2 _24091_ (.A0(\w[19][6] ),
    .A1(\w[17][6] ),
    .A2(\w[23][6] ),
    .A3(\w[21][6] ),
    .S0(net359),
    .S1(net309),
    .X(_09972_));
 sky130_fd_sc_hd__mux4_2 _24092_ (.A0(\w[27][6] ),
    .A1(\w[25][6] ),
    .A2(\w[31][6] ),
    .A3(\w[29][6] ),
    .S0(net359),
    .S1(net309),
    .X(_09973_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_551 ();
 sky130_fd_sc_hd__mux4_2 _24094_ (.A0(\w[3][6] ),
    .A1(\w[1][6] ),
    .A2(\w[7][6] ),
    .A3(\w[5][6] ),
    .S0(net359),
    .S1(net309),
    .X(_09975_));
 sky130_fd_sc_hd__mux4_2 _24095_ (.A0(\w[11][6] ),
    .A1(\w[9][6] ),
    .A2(\w[15][6] ),
    .A3(\w[13][6] ),
    .S0(net359),
    .S1(net309),
    .X(_09976_));
 sky130_fd_sc_hd__mux4_2 _24096_ (.A0(_09972_),
    .A1(_09973_),
    .A2(_09975_),
    .A3(_09976_),
    .S0(net333),
    .S1(net327),
    .X(_09977_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_550 ();
 sky130_fd_sc_hd__mux4_2 _24098_ (.A0(\w[51][6] ),
    .A1(\w[49][6] ),
    .A2(\w[55][6] ),
    .A3(\w[53][6] ),
    .S0(net362),
    .S1(net310),
    .X(_09979_));
 sky130_fd_sc_hd__mux4_2 _24099_ (.A0(\w[59][6] ),
    .A1(\w[57][6] ),
    .A2(\w[63][6] ),
    .A3(\w[61][6] ),
    .S0(net362),
    .S1(net310),
    .X(_09980_));
 sky130_fd_sc_hd__mux4_2 _24100_ (.A0(\w[35][6] ),
    .A1(\w[33][6] ),
    .A2(\w[39][6] ),
    .A3(\w[37][6] ),
    .S0(net362),
    .S1(net310),
    .X(_09981_));
 sky130_fd_sc_hd__mux4_2 _24101_ (.A0(\w[43][6] ),
    .A1(\w[41][6] ),
    .A2(\w[47][6] ),
    .A3(\w[45][6] ),
    .S0(net362),
    .S1(net310),
    .X(_09982_));
 sky130_fd_sc_hd__mux4_2 _24102_ (.A0(_09979_),
    .A1(_09980_),
    .A2(_09981_),
    .A3(_09982_),
    .S0(net336),
    .S1(net328),
    .X(_09983_));
 sky130_fd_sc_hd__mux2i_1 _24103_ (.A0(_09977_),
    .A1(_09983_),
    .S(net292),
    .Y(_09984_));
 sky130_fd_sc_hd__nand2_2 _24104_ (.A(net347),
    .B(\w[1][6] ),
    .Y(_09985_));
 sky130_fd_sc_hd__o21ai_4 _24105_ (.A1(net285),
    .A2(_09984_),
    .B1(_09985_),
    .Y(_00060_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_549 ();
 sky130_fd_sc_hd__mux4_2 _24107_ (.A0(\w[19][7] ),
    .A1(\w[17][7] ),
    .A2(\w[23][7] ),
    .A3(\w[21][7] ),
    .S0(net360),
    .S1(net308),
    .X(_09987_));
 sky130_fd_sc_hd__mux4_2 _24108_ (.A0(\w[27][7] ),
    .A1(\w[25][7] ),
    .A2(\w[31][7] ),
    .A3(\w[29][7] ),
    .S0(net360),
    .S1(net308),
    .X(_09988_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_548 ();
 sky130_fd_sc_hd__mux4_2 _24110_ (.A0(\w[3][7] ),
    .A1(\w[1][7] ),
    .A2(\w[7][7] ),
    .A3(\w[5][7] ),
    .S0(net360),
    .S1(net308),
    .X(_09990_));
 sky130_fd_sc_hd__mux4_2 _24111_ (.A0(\w[11][7] ),
    .A1(\w[9][7] ),
    .A2(\w[15][7] ),
    .A3(\w[13][7] ),
    .S0(net360),
    .S1(net308),
    .X(_09991_));
 sky130_fd_sc_hd__mux4_2 _24112_ (.A0(_09987_),
    .A1(_09988_),
    .A2(_09990_),
    .A3(_09991_),
    .S0(net335),
    .S1(net330),
    .X(_09992_));
 sky130_fd_sc_hd__mux4_2 _24113_ (.A0(\w[51][7] ),
    .A1(\w[49][7] ),
    .A2(\w[55][7] ),
    .A3(\w[53][7] ),
    .S0(net360),
    .S1(net308),
    .X(_09993_));
 sky130_fd_sc_hd__mux4_2 _24114_ (.A0(\w[59][7] ),
    .A1(\w[57][7] ),
    .A2(\w[63][7] ),
    .A3(\w[61][7] ),
    .S0(net360),
    .S1(net308),
    .X(_09994_));
 sky130_fd_sc_hd__mux4_2 _24115_ (.A0(\w[35][7] ),
    .A1(\w[33][7] ),
    .A2(\w[39][7] ),
    .A3(\w[37][7] ),
    .S0(net360),
    .S1(net308),
    .X(_09995_));
 sky130_fd_sc_hd__mux4_2 _24116_ (.A0(\w[43][7] ),
    .A1(\w[41][7] ),
    .A2(\w[47][7] ),
    .A3(\w[45][7] ),
    .S0(net360),
    .S1(net308),
    .X(_09996_));
 sky130_fd_sc_hd__mux4_2 _24117_ (.A0(_09993_),
    .A1(_09994_),
    .A2(_09995_),
    .A3(_09996_),
    .S0(net335),
    .S1(net330),
    .X(_09997_));
 sky130_fd_sc_hd__mux2i_1 _24118_ (.A0(_09992_),
    .A1(_09997_),
    .S(net295),
    .Y(_09998_));
 sky130_fd_sc_hd__nand2_2 _24119_ (.A(net347),
    .B(\w[1][7] ),
    .Y(_09999_));
 sky130_fd_sc_hd__o21ai_4 _24120_ (.A1(net285),
    .A2(_09998_),
    .B1(_09999_),
    .Y(_00061_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_547 ();
 sky130_fd_sc_hd__mux4_2 _24122_ (.A0(\w[19][8] ),
    .A1(\w[17][8] ),
    .A2(\w[23][8] ),
    .A3(\w[21][8] ),
    .S0(net363),
    .S1(net311),
    .X(_10001_));
 sky130_fd_sc_hd__mux4_2 _24123_ (.A0(\w[27][8] ),
    .A1(\w[25][8] ),
    .A2(\w[31][8] ),
    .A3(\w[29][8] ),
    .S0(net363),
    .S1(net311),
    .X(_10002_));
 sky130_fd_sc_hd__mux4_2 _24124_ (.A0(\w[3][8] ),
    .A1(\w[1][8] ),
    .A2(\w[7][8] ),
    .A3(\w[5][8] ),
    .S0(net363),
    .S1(net311),
    .X(_10003_));
 sky130_fd_sc_hd__mux4_2 _24125_ (.A0(\w[11][8] ),
    .A1(\w[9][8] ),
    .A2(\w[15][8] ),
    .A3(\w[13][8] ),
    .S0(net363),
    .S1(net311),
    .X(_10004_));
 sky130_fd_sc_hd__mux4_2 _24126_ (.A0(_10001_),
    .A1(_10002_),
    .A2(_10003_),
    .A3(_10004_),
    .S0(net334),
    .S1(net327),
    .X(_10005_));
 sky130_fd_sc_hd__mux4_2 _24127_ (.A0(\w[51][8] ),
    .A1(\w[49][8] ),
    .A2(\w[55][8] ),
    .A3(\w[53][8] ),
    .S0(net362),
    .S1(net309),
    .X(_10006_));
 sky130_fd_sc_hd__mux4_2 _24128_ (.A0(\w[59][8] ),
    .A1(\w[57][8] ),
    .A2(\w[63][8] ),
    .A3(\w[61][8] ),
    .S0(net362),
    .S1(net309),
    .X(_10007_));
 sky130_fd_sc_hd__mux4_2 _24129_ (.A0(\w[35][8] ),
    .A1(\w[33][8] ),
    .A2(\w[39][8] ),
    .A3(\w[37][8] ),
    .S0(net359),
    .S1(net309),
    .X(_10008_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_546 ();
 sky130_fd_sc_hd__mux4_2 _24131_ (.A0(\w[43][8] ),
    .A1(\w[41][8] ),
    .A2(\w[47][8] ),
    .A3(\w[45][8] ),
    .S0(net362),
    .S1(net309),
    .X(_10010_));
 sky130_fd_sc_hd__mux4_2 _24132_ (.A0(_10006_),
    .A1(_10007_),
    .A2(_10008_),
    .A3(_10010_),
    .S0(net334),
    .S1(net328),
    .X(_10011_));
 sky130_fd_sc_hd__mux2i_1 _24133_ (.A0(_10005_),
    .A1(_10011_),
    .S(net292),
    .Y(_10012_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_544 ();
 sky130_fd_sc_hd__nand2_2 _24136_ (.A(net347),
    .B(\w[1][8] ),
    .Y(_10015_));
 sky130_fd_sc_hd__o21ai_4 _24137_ (.A1(net285),
    .A2(_10012_),
    .B1(_10015_),
    .Y(_00062_));
 sky130_fd_sc_hd__mux4_2 _24138_ (.A0(\w[19][9] ),
    .A1(\w[17][9] ),
    .A2(\w[23][9] ),
    .A3(\w[21][9] ),
    .S0(net364),
    .S1(net312),
    .X(_10016_));
 sky130_fd_sc_hd__mux4_2 _24139_ (.A0(\w[27][9] ),
    .A1(\w[25][9] ),
    .A2(\w[31][9] ),
    .A3(\w[29][9] ),
    .S0(net364),
    .S1(net312),
    .X(_10017_));
 sky130_fd_sc_hd__mux4_2 _24140_ (.A0(\w[3][9] ),
    .A1(\w[1][9] ),
    .A2(\w[7][9] ),
    .A3(\w[5][9] ),
    .S0(net364),
    .S1(net312),
    .X(_10018_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_543 ();
 sky130_fd_sc_hd__mux4_2 _24142_ (.A0(\w[11][9] ),
    .A1(\w[9][9] ),
    .A2(\w[15][9] ),
    .A3(\w[13][9] ),
    .S0(net364),
    .S1(net312),
    .X(_10020_));
 sky130_fd_sc_hd__mux4_2 _24143_ (.A0(_10016_),
    .A1(_10017_),
    .A2(_10018_),
    .A3(_10020_),
    .S0(net332),
    .S1(net330),
    .X(_10021_));
 sky130_fd_sc_hd__mux4_2 _24144_ (.A0(\w[51][9] ),
    .A1(\w[49][9] ),
    .A2(\w[55][9] ),
    .A3(\w[53][9] ),
    .S0(net364),
    .S1(net308),
    .X(_10022_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_542 ();
 sky130_fd_sc_hd__mux4_2 _24146_ (.A0(\w[59][9] ),
    .A1(\w[57][9] ),
    .A2(\w[63][9] ),
    .A3(\w[61][9] ),
    .S0(net364),
    .S1(net308),
    .X(_10024_));
 sky130_fd_sc_hd__mux4_2 _24147_ (.A0(\w[35][9] ),
    .A1(\w[33][9] ),
    .A2(\w[39][9] ),
    .A3(\w[37][9] ),
    .S0(net364),
    .S1(net308),
    .X(_10025_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_541 ();
 sky130_fd_sc_hd__mux4_2 _24149_ (.A0(\w[43][9] ),
    .A1(\w[41][9] ),
    .A2(\w[47][9] ),
    .A3(\w[45][9] ),
    .S0(net364),
    .S1(net308),
    .X(_10027_));
 sky130_fd_sc_hd__mux4_2 _24150_ (.A0(_10022_),
    .A1(_10024_),
    .A2(_10025_),
    .A3(_10027_),
    .S0(net335),
    .S1(net330),
    .X(_10028_));
 sky130_fd_sc_hd__mux2i_1 _24151_ (.A0(_10021_),
    .A1(_10028_),
    .S(net295),
    .Y(_10029_));
 sky130_fd_sc_hd__nand2_2 _24152_ (.A(net347),
    .B(\w[1][9] ),
    .Y(_10030_));
 sky130_fd_sc_hd__o21ai_4 _24153_ (.A1(net287),
    .A2(_10029_),
    .B1(_10030_),
    .Y(_00063_));
 sky130_fd_sc_hd__mux4_2 _24154_ (.A0(\w[19][10] ),
    .A1(\w[17][10] ),
    .A2(\w[23][10] ),
    .A3(\w[21][10] ),
    .S0(net361),
    .S1(net311),
    .X(_10031_));
 sky130_fd_sc_hd__mux4_2 _24155_ (.A0(\w[27][10] ),
    .A1(\w[25][10] ),
    .A2(\w[31][10] ),
    .A3(\w[29][10] ),
    .S0(net361),
    .S1(net311),
    .X(_10032_));
 sky130_fd_sc_hd__mux4_2 _24156_ (.A0(\w[3][10] ),
    .A1(\w[1][10] ),
    .A2(\w[7][10] ),
    .A3(\w[5][10] ),
    .S0(net361),
    .S1(net311),
    .X(_10033_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_540 ();
 sky130_fd_sc_hd__mux4_2 _24158_ (.A0(\w[11][10] ),
    .A1(\w[9][10] ),
    .A2(\w[15][10] ),
    .A3(\w[13][10] ),
    .S0(net361),
    .S1(net311),
    .X(_10035_));
 sky130_fd_sc_hd__mux4_2 _24159_ (.A0(_10031_),
    .A1(_10032_),
    .A2(_10033_),
    .A3(_10035_),
    .S0(net337),
    .S1(net329),
    .X(_10036_));
 sky130_fd_sc_hd__mux4_2 _24160_ (.A0(\w[51][10] ),
    .A1(\w[49][10] ),
    .A2(\w[55][10] ),
    .A3(\w[53][10] ),
    .S0(net362),
    .S1(net310),
    .X(_10037_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_539 ();
 sky130_fd_sc_hd__mux4_2 _24162_ (.A0(\w[59][10] ),
    .A1(\w[57][10] ),
    .A2(\w[63][10] ),
    .A3(\w[61][10] ),
    .S0(net362),
    .S1(net310),
    .X(_10039_));
 sky130_fd_sc_hd__mux4_2 _24163_ (.A0(\w[35][10] ),
    .A1(\w[33][10] ),
    .A2(\w[39][10] ),
    .A3(\w[37][10] ),
    .S0(net362),
    .S1(net310),
    .X(_10040_));
 sky130_fd_sc_hd__mux4_2 _24164_ (.A0(\w[43][10] ),
    .A1(\w[41][10] ),
    .A2(\w[47][10] ),
    .A3(\w[45][10] ),
    .S0(net362),
    .S1(net310),
    .X(_10041_));
 sky130_fd_sc_hd__mux4_2 _24165_ (.A0(_10037_),
    .A1(_10039_),
    .A2(_10040_),
    .A3(_10041_),
    .S0(net336),
    .S1(net328),
    .X(_10042_));
 sky130_fd_sc_hd__mux2i_1 _24166_ (.A0(_10036_),
    .A1(_10042_),
    .S(net293),
    .Y(_10043_));
 sky130_fd_sc_hd__nand2_1 _24167_ (.A(net347),
    .B(\w[1][10] ),
    .Y(_10044_));
 sky130_fd_sc_hd__o21ai_0 _24168_ (.A1(net285),
    .A2(_10043_),
    .B1(_10044_),
    .Y(_00033_));
 sky130_fd_sc_hd__mux4_2 _24169_ (.A0(\w[19][11] ),
    .A1(\w[17][11] ),
    .A2(\w[23][11] ),
    .A3(\w[21][11] ),
    .S0(net363),
    .S1(net311),
    .X(_10045_));
 sky130_fd_sc_hd__mux4_2 _24170_ (.A0(\w[27][11] ),
    .A1(\w[25][11] ),
    .A2(\w[31][11] ),
    .A3(\w[29][11] ),
    .S0(net363),
    .S1(net311),
    .X(_10046_));
 sky130_fd_sc_hd__mux4_2 _24171_ (.A0(\w[3][11] ),
    .A1(\w[1][11] ),
    .A2(\w[7][11] ),
    .A3(\w[5][11] ),
    .S0(net363),
    .S1(net311),
    .X(_10047_));
 sky130_fd_sc_hd__mux4_2 _24172_ (.A0(\w[11][11] ),
    .A1(\w[9][11] ),
    .A2(\w[15][11] ),
    .A3(\w[13][11] ),
    .S0(net363),
    .S1(net311),
    .X(_10048_));
 sky130_fd_sc_hd__mux4_2 _24173_ (.A0(_10045_),
    .A1(_10046_),
    .A2(_10047_),
    .A3(_10048_),
    .S0(net334),
    .S1(net329),
    .X(_10049_));
 sky130_fd_sc_hd__mux4_2 _24174_ (.A0(\w[51][11] ),
    .A1(\w[49][11] ),
    .A2(\w[55][11] ),
    .A3(\w[53][11] ),
    .S0(net364),
    .S1(net312),
    .X(_10050_));
 sky130_fd_sc_hd__mux4_2 _24175_ (.A0(\w[59][11] ),
    .A1(\w[57][11] ),
    .A2(\w[63][11] ),
    .A3(\w[61][11] ),
    .S0(net364),
    .S1(net312),
    .X(_10051_));
 sky130_fd_sc_hd__mux4_2 _24176_ (.A0(\w[35][11] ),
    .A1(\w[33][11] ),
    .A2(\w[39][11] ),
    .A3(\w[37][11] ),
    .S0(net364),
    .S1(net312),
    .X(_10052_));
 sky130_fd_sc_hd__mux4_2 _24177_ (.A0(\w[43][11] ),
    .A1(\w[41][11] ),
    .A2(\w[47][11] ),
    .A3(\w[45][11] ),
    .S0(net364),
    .S1(net312),
    .X(_10053_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_538 ();
 sky130_fd_sc_hd__mux4_2 _24179_ (.A0(_10050_),
    .A1(_10051_),
    .A2(_10052_),
    .A3(_10053_),
    .S0(_09854_),
    .S1(net331),
    .X(_10055_));
 sky130_fd_sc_hd__mux2i_1 _24180_ (.A0(_10049_),
    .A1(_10055_),
    .S(net292),
    .Y(_10056_));
 sky130_fd_sc_hd__nand2_2 _24181_ (.A(net347),
    .B(\w[1][11] ),
    .Y(_10057_));
 sky130_fd_sc_hd__o21ai_4 _24182_ (.A1(net285),
    .A2(_10056_),
    .B1(_10057_),
    .Y(_00034_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_537 ();
 sky130_fd_sc_hd__mux4_2 _24184_ (.A0(\w[19][12] ),
    .A1(\w[17][12] ),
    .A2(\w[23][12] ),
    .A3(\w[21][12] ),
    .S0(net363),
    .S1(net311),
    .X(_10059_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_536 ();
 sky130_fd_sc_hd__mux4_2 _24186_ (.A0(\w[27][12] ),
    .A1(\w[25][12] ),
    .A2(\w[31][12] ),
    .A3(\w[29][12] ),
    .S0(net363),
    .S1(net311),
    .X(_10061_));
 sky130_fd_sc_hd__mux4_2 _24187_ (.A0(\w[3][12] ),
    .A1(\w[1][12] ),
    .A2(\w[7][12] ),
    .A3(\w[5][12] ),
    .S0(net363),
    .S1(net311),
    .X(_10062_));
 sky130_fd_sc_hd__mux4_2 _24188_ (.A0(\w[11][12] ),
    .A1(\w[9][12] ),
    .A2(\w[15][12] ),
    .A3(\w[13][12] ),
    .S0(net363),
    .S1(net311),
    .X(_10063_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_535 ();
 sky130_fd_sc_hd__mux4_2 _24190_ (.A0(_10059_),
    .A1(_10061_),
    .A2(_10062_),
    .A3(_10063_),
    .S0(net334),
    .S1(net327),
    .X(_10065_));
 sky130_fd_sc_hd__mux4_2 _24191_ (.A0(\w[51][12] ),
    .A1(\w[49][12] ),
    .A2(\w[55][12] ),
    .A3(\w[53][12] ),
    .S0(net360),
    .S1(_00657_),
    .X(_10066_));
 sky130_fd_sc_hd__mux4_2 _24192_ (.A0(\w[59][12] ),
    .A1(\w[57][12] ),
    .A2(\w[63][12] ),
    .A3(\w[61][12] ),
    .S0(net360),
    .S1(_00657_),
    .X(_10067_));
 sky130_fd_sc_hd__mux4_2 _24193_ (.A0(\w[35][12] ),
    .A1(\w[33][12] ),
    .A2(\w[39][12] ),
    .A3(\w[37][12] ),
    .S0(net362),
    .S1(_00657_),
    .X(_10068_));
 sky130_fd_sc_hd__mux4_2 _24194_ (.A0(\w[43][12] ),
    .A1(\w[41][12] ),
    .A2(\w[47][12] ),
    .A3(\w[45][12] ),
    .S0(net362),
    .S1(net310),
    .X(_10069_));
 sky130_fd_sc_hd__mux4_2 _24195_ (.A0(_10066_),
    .A1(_10067_),
    .A2(_10068_),
    .A3(_10069_),
    .S0(net338),
    .S1(_09857_),
    .X(_10070_));
 sky130_fd_sc_hd__mux2i_1 _24196_ (.A0(_10065_),
    .A1(_10070_),
    .S(net292),
    .Y(_10071_));
 sky130_fd_sc_hd__nand2_2 _24197_ (.A(net347),
    .B(\w[1][12] ),
    .Y(_10072_));
 sky130_fd_sc_hd__o21ai_4 _24198_ (.A1(net285),
    .A2(_10071_),
    .B1(_10072_),
    .Y(_00035_));
 sky130_fd_sc_hd__mux4_2 _24199_ (.A0(\w[19][13] ),
    .A1(\w[17][13] ),
    .A2(\w[23][13] ),
    .A3(\w[21][13] ),
    .S0(net361),
    .S1(net311),
    .X(_10073_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_534 ();
 sky130_fd_sc_hd__mux4_2 _24201_ (.A0(\w[27][13] ),
    .A1(\w[25][13] ),
    .A2(\w[31][13] ),
    .A3(\w[29][13] ),
    .S0(net361),
    .S1(net311),
    .X(_10075_));
 sky130_fd_sc_hd__mux4_2 _24202_ (.A0(\w[3][13] ),
    .A1(\w[1][13] ),
    .A2(\w[7][13] ),
    .A3(\w[5][13] ),
    .S0(net361),
    .S1(net311),
    .X(_10076_));
 sky130_fd_sc_hd__mux4_2 _24203_ (.A0(\w[11][13] ),
    .A1(\w[9][13] ),
    .A2(\w[15][13] ),
    .A3(\w[13][13] ),
    .S0(net361),
    .S1(net311),
    .X(_10077_));
 sky130_fd_sc_hd__mux4_2 _24204_ (.A0(_10073_),
    .A1(_10075_),
    .A2(_10076_),
    .A3(_10077_),
    .S0(net337),
    .S1(net329),
    .X(_10078_));
 sky130_fd_sc_hd__mux4_2 _24205_ (.A0(\w[51][13] ),
    .A1(\w[49][13] ),
    .A2(\w[55][13] ),
    .A3(\w[53][13] ),
    .S0(net363),
    .S1(_00657_),
    .X(_10079_));
 sky130_fd_sc_hd__mux4_2 _24206_ (.A0(\w[59][13] ),
    .A1(\w[57][13] ),
    .A2(\w[63][13] ),
    .A3(\w[61][13] ),
    .S0(net363),
    .S1(_00657_),
    .X(_10080_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_533 ();
 sky130_fd_sc_hd__mux4_2 _24208_ (.A0(\w[35][13] ),
    .A1(\w[33][13] ),
    .A2(\w[39][13] ),
    .A3(\w[37][13] ),
    .S0(net363),
    .S1(_00657_),
    .X(_10082_));
 sky130_fd_sc_hd__mux4_2 _24209_ (.A0(\w[43][13] ),
    .A1(\w[41][13] ),
    .A2(\w[47][13] ),
    .A3(\w[45][13] ),
    .S0(net363),
    .S1(_00657_),
    .X(_10083_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_532 ();
 sky130_fd_sc_hd__mux4_2 _24211_ (.A0(_10079_),
    .A1(_10080_),
    .A2(_10082_),
    .A3(_10083_),
    .S0(_09854_),
    .S1(_09857_),
    .X(_10085_));
 sky130_fd_sc_hd__mux2i_1 _24212_ (.A0(_10078_),
    .A1(_10085_),
    .S(net293),
    .Y(_10086_));
 sky130_fd_sc_hd__nand2_1 _24213_ (.A(net347),
    .B(\w[1][13] ),
    .Y(_10087_));
 sky130_fd_sc_hd__o21ai_0 _24214_ (.A1(net285),
    .A2(_10086_),
    .B1(_10087_),
    .Y(_00036_));
 sky130_fd_sc_hd__mux4_2 _24215_ (.A0(\w[19][14] ),
    .A1(\w[17][14] ),
    .A2(\w[23][14] ),
    .A3(\w[21][14] ),
    .S0(net359),
    .S1(net309),
    .X(_10088_));
 sky130_fd_sc_hd__mux4_2 _24216_ (.A0(\w[27][14] ),
    .A1(\w[25][14] ),
    .A2(\w[31][14] ),
    .A3(\w[29][14] ),
    .S0(net359),
    .S1(net309),
    .X(_10089_));
 sky130_fd_sc_hd__mux4_2 _24217_ (.A0(\w[3][14] ),
    .A1(\w[1][14] ),
    .A2(\w[7][14] ),
    .A3(\w[5][14] ),
    .S0(net359),
    .S1(net309),
    .X(_10090_));
 sky130_fd_sc_hd__mux4_2 _24218_ (.A0(\w[11][14] ),
    .A1(\w[9][14] ),
    .A2(\w[15][14] ),
    .A3(\w[13][14] ),
    .S0(net359),
    .S1(net309),
    .X(_10091_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_531 ();
 sky130_fd_sc_hd__mux4_2 _24220_ (.A0(_10088_),
    .A1(_10089_),
    .A2(_10090_),
    .A3(_10091_),
    .S0(net334),
    .S1(net327),
    .X(_10093_));
 sky130_fd_sc_hd__mux4_2 _24221_ (.A0(\w[51][14] ),
    .A1(\w[49][14] ),
    .A2(\w[55][14] ),
    .A3(\w[53][14] ),
    .S0(net362),
    .S1(net309),
    .X(_10094_));
 sky130_fd_sc_hd__mux4_2 _24222_ (.A0(\w[59][14] ),
    .A1(\w[57][14] ),
    .A2(\w[63][14] ),
    .A3(\w[61][14] ),
    .S0(net362),
    .S1(net309),
    .X(_10095_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_530 ();
 sky130_fd_sc_hd__mux4_2 _24224_ (.A0(\w[35][14] ),
    .A1(\w[33][14] ),
    .A2(\w[39][14] ),
    .A3(\w[37][14] ),
    .S0(net362),
    .S1(net309),
    .X(_10097_));
 sky130_fd_sc_hd__mux4_2 _24225_ (.A0(\w[43][14] ),
    .A1(\w[41][14] ),
    .A2(\w[47][14] ),
    .A3(\w[45][14] ),
    .S0(net362),
    .S1(net309),
    .X(_10098_));
 sky130_fd_sc_hd__mux4_2 _24226_ (.A0(_10094_),
    .A1(_10095_),
    .A2(_10097_),
    .A3(_10098_),
    .S0(net336),
    .S1(net326),
    .X(_10099_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_529 ();
 sky130_fd_sc_hd__mux2i_1 _24228_ (.A0(_10093_),
    .A1(_10099_),
    .S(net292),
    .Y(_10101_));
 sky130_fd_sc_hd__nand2_2 _24229_ (.A(net347),
    .B(\w[1][14] ),
    .Y(_10102_));
 sky130_fd_sc_hd__o21ai_4 _24230_ (.A1(net285),
    .A2(_10101_),
    .B1(_10102_),
    .Y(_00037_));
 sky130_fd_sc_hd__mux4_2 _24231_ (.A0(\w[19][15] ),
    .A1(\w[17][15] ),
    .A2(\w[23][15] ),
    .A3(\w[21][15] ),
    .S0(net357),
    .S1(net312),
    .X(_10103_));
 sky130_fd_sc_hd__mux4_2 _24232_ (.A0(\w[27][15] ),
    .A1(\w[25][15] ),
    .A2(\w[31][15] ),
    .A3(\w[29][15] ),
    .S0(net357),
    .S1(net312),
    .X(_10104_));
 sky130_fd_sc_hd__mux4_2 _24233_ (.A0(\w[3][15] ),
    .A1(\w[1][15] ),
    .A2(\w[7][15] ),
    .A3(\w[5][15] ),
    .S0(net357),
    .S1(net312),
    .X(_10105_));
 sky130_fd_sc_hd__mux4_2 _24234_ (.A0(\w[11][15] ),
    .A1(\w[9][15] ),
    .A2(\w[15][15] ),
    .A3(\w[13][15] ),
    .S0(net357),
    .S1(net312),
    .X(_10106_));
 sky130_fd_sc_hd__mux4_2 _24235_ (.A0(_10103_),
    .A1(_10104_),
    .A2(_10105_),
    .A3(_10106_),
    .S0(net332),
    .S1(net331),
    .X(_10107_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_528 ();
 sky130_fd_sc_hd__mux4_2 _24237_ (.A0(\w[51][15] ),
    .A1(\w[49][15] ),
    .A2(\w[55][15] ),
    .A3(\w[53][15] ),
    .S0(net357),
    .S1(net312),
    .X(_10109_));
 sky130_fd_sc_hd__mux4_2 _24238_ (.A0(\w[59][15] ),
    .A1(\w[57][15] ),
    .A2(\w[63][15] ),
    .A3(\w[61][15] ),
    .S0(net357),
    .S1(net312),
    .X(_10110_));
 sky130_fd_sc_hd__mux4_2 _24239_ (.A0(\w[35][15] ),
    .A1(\w[33][15] ),
    .A2(\w[39][15] ),
    .A3(\w[37][15] ),
    .S0(net357),
    .S1(net312),
    .X(_10111_));
 sky130_fd_sc_hd__mux4_2 _24240_ (.A0(\w[43][15] ),
    .A1(\w[41][15] ),
    .A2(\w[47][15] ),
    .A3(\w[45][15] ),
    .S0(net357),
    .S1(net312),
    .X(_10112_));
 sky130_fd_sc_hd__mux4_2 _24241_ (.A0(_10109_),
    .A1(_10110_),
    .A2(_10111_),
    .A3(_10112_),
    .S0(net332),
    .S1(net331),
    .X(_10113_));
 sky130_fd_sc_hd__mux2i_1 _24242_ (.A0(_10107_),
    .A1(_10113_),
    .S(net295),
    .Y(_10114_));
 sky130_fd_sc_hd__nand2_2 _24243_ (.A(net349),
    .B(\w[1][15] ),
    .Y(_10115_));
 sky130_fd_sc_hd__o21ai_4 _24244_ (.A1(net287),
    .A2(_10114_),
    .B1(_10115_),
    .Y(_00038_));
 sky130_fd_sc_hd__mux4_2 _24245_ (.A0(\w[19][16] ),
    .A1(\w[17][16] ),
    .A2(\w[23][16] ),
    .A3(\w[21][16] ),
    .S0(net359),
    .S1(net309),
    .X(_10116_));
 sky130_fd_sc_hd__mux4_2 _24246_ (.A0(\w[27][16] ),
    .A1(\w[25][16] ),
    .A2(\w[31][16] ),
    .A3(\w[29][16] ),
    .S0(net359),
    .S1(net309),
    .X(_10117_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_527 ();
 sky130_fd_sc_hd__mux4_2 _24248_ (.A0(\w[3][16] ),
    .A1(\w[1][16] ),
    .A2(\w[7][16] ),
    .A3(\w[5][16] ),
    .S0(net359),
    .S1(net309),
    .X(_10119_));
 sky130_fd_sc_hd__mux4_2 _24249_ (.A0(\w[11][16] ),
    .A1(\w[9][16] ),
    .A2(\w[15][16] ),
    .A3(\w[13][16] ),
    .S0(net359),
    .S1(net309),
    .X(_10120_));
 sky130_fd_sc_hd__mux4_2 _24250_ (.A0(_10116_),
    .A1(_10117_),
    .A2(_10119_),
    .A3(_10120_),
    .S0(net333),
    .S1(net327),
    .X(_10121_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_526 ();
 sky130_fd_sc_hd__mux4_2 _24252_ (.A0(\w[51][16] ),
    .A1(\w[49][16] ),
    .A2(\w[55][16] ),
    .A3(\w[53][16] ),
    .S0(net360),
    .S1(net308),
    .X(_10123_));
 sky130_fd_sc_hd__mux4_2 _24253_ (.A0(\w[59][16] ),
    .A1(\w[57][16] ),
    .A2(\w[63][16] ),
    .A3(\w[61][16] ),
    .S0(net360),
    .S1(net308),
    .X(_10124_));
 sky130_fd_sc_hd__mux4_2 _24254_ (.A0(\w[35][16] ),
    .A1(\w[33][16] ),
    .A2(\w[39][16] ),
    .A3(\w[37][16] ),
    .S0(net360),
    .S1(_00657_),
    .X(_10125_));
 sky130_fd_sc_hd__mux4_2 _24255_ (.A0(\w[43][16] ),
    .A1(\w[41][16] ),
    .A2(\w[47][16] ),
    .A3(\w[45][16] ),
    .S0(net360),
    .S1(net308),
    .X(_10126_));
 sky130_fd_sc_hd__mux4_2 _24256_ (.A0(_10123_),
    .A1(_10124_),
    .A2(_10125_),
    .A3(_10126_),
    .S0(net335),
    .S1(net328),
    .X(_10127_));
 sky130_fd_sc_hd__mux2i_1 _24257_ (.A0(_10121_),
    .A1(_10127_),
    .S(net292),
    .Y(_10128_));
 sky130_fd_sc_hd__nand2_2 _24258_ (.A(net347),
    .B(\w[1][16] ),
    .Y(_10129_));
 sky130_fd_sc_hd__o21ai_4 _24259_ (.A1(net285),
    .A2(_10128_),
    .B1(_10129_),
    .Y(_00039_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_525 ();
 sky130_fd_sc_hd__mux4_2 _24261_ (.A0(\w[19][17] ),
    .A1(\w[17][17] ),
    .A2(\w[23][17] ),
    .A3(\w[21][17] ),
    .S0(net359),
    .S1(net309),
    .X(_10131_));
 sky130_fd_sc_hd__mux4_2 _24262_ (.A0(\w[27][17] ),
    .A1(\w[25][17] ),
    .A2(\w[31][17] ),
    .A3(\w[29][17] ),
    .S0(net359),
    .S1(net309),
    .X(_10132_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_524 ();
 sky130_fd_sc_hd__mux4_2 _24264_ (.A0(\w[3][17] ),
    .A1(\w[1][17] ),
    .A2(\w[7][17] ),
    .A3(\w[5][17] ),
    .S0(net359),
    .S1(net309),
    .X(_10134_));
 sky130_fd_sc_hd__mux4_2 _24265_ (.A0(\w[11][17] ),
    .A1(\w[9][17] ),
    .A2(\w[15][17] ),
    .A3(\w[13][17] ),
    .S0(net359),
    .S1(net309),
    .X(_10135_));
 sky130_fd_sc_hd__mux4_2 _24266_ (.A0(_10131_),
    .A1(_10132_),
    .A2(_10134_),
    .A3(_10135_),
    .S0(net333),
    .S1(net327),
    .X(_10136_));
 sky130_fd_sc_hd__mux4_2 _24267_ (.A0(\w[51][17] ),
    .A1(\w[49][17] ),
    .A2(\w[55][17] ),
    .A3(\w[53][17] ),
    .S0(net358),
    .S1(net310),
    .X(_10137_));
 sky130_fd_sc_hd__mux4_2 _24268_ (.A0(\w[59][17] ),
    .A1(\w[57][17] ),
    .A2(\w[63][17] ),
    .A3(\w[61][17] ),
    .S0(net358),
    .S1(net310),
    .X(_10138_));
 sky130_fd_sc_hd__mux4_2 _24269_ (.A0(\w[35][17] ),
    .A1(\w[33][17] ),
    .A2(\w[39][17] ),
    .A3(\w[37][17] ),
    .S0(net358),
    .S1(net310),
    .X(_10139_));
 sky130_fd_sc_hd__mux4_2 _24270_ (.A0(\w[43][17] ),
    .A1(\w[41][17] ),
    .A2(\w[47][17] ),
    .A3(\w[45][17] ),
    .S0(net358),
    .S1(net310),
    .X(_10140_));
 sky130_fd_sc_hd__mux4_2 _24271_ (.A0(_10137_),
    .A1(_10138_),
    .A2(_10139_),
    .A3(_10140_),
    .S0(net336),
    .S1(net326),
    .X(_10141_));
 sky130_fd_sc_hd__mux2i_1 _24272_ (.A0(_10136_),
    .A1(_10141_),
    .S(net292),
    .Y(_10142_));
 sky130_fd_sc_hd__nand2_2 _24273_ (.A(net347),
    .B(\w[1][17] ),
    .Y(_10143_));
 sky130_fd_sc_hd__o21ai_4 _24274_ (.A1(net285),
    .A2(_10142_),
    .B1(_10143_),
    .Y(_00040_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_523 ();
 sky130_fd_sc_hd__mux4_2 _24276_ (.A0(\w[19][18] ),
    .A1(\w[17][18] ),
    .A2(\w[23][18] ),
    .A3(\w[21][18] ),
    .S0(net361),
    .S1(net311),
    .X(_10145_));
 sky130_fd_sc_hd__mux4_2 _24277_ (.A0(\w[27][18] ),
    .A1(\w[25][18] ),
    .A2(\w[31][18] ),
    .A3(\w[29][18] ),
    .S0(net361),
    .S1(net311),
    .X(_10146_));
 sky130_fd_sc_hd__mux4_2 _24278_ (.A0(\w[3][18] ),
    .A1(\w[1][18] ),
    .A2(\w[7][18] ),
    .A3(\w[5][18] ),
    .S0(net361),
    .S1(net311),
    .X(_10147_));
 sky130_fd_sc_hd__mux4_2 _24279_ (.A0(\w[11][18] ),
    .A1(\w[9][18] ),
    .A2(\w[15][18] ),
    .A3(\w[13][18] ),
    .S0(net361),
    .S1(net311),
    .X(_10148_));
 sky130_fd_sc_hd__mux4_2 _24280_ (.A0(_10145_),
    .A1(_10146_),
    .A2(_10147_),
    .A3(_10148_),
    .S0(net337),
    .S1(net329),
    .X(_10149_));
 sky130_fd_sc_hd__mux4_2 _24281_ (.A0(\w[51][18] ),
    .A1(\w[49][18] ),
    .A2(\w[55][18] ),
    .A3(\w[53][18] ),
    .S0(net363),
    .S1(net311),
    .X(_10150_));
 sky130_fd_sc_hd__mux4_2 _24282_ (.A0(\w[59][18] ),
    .A1(\w[57][18] ),
    .A2(\w[63][18] ),
    .A3(\w[61][18] ),
    .S0(net363),
    .S1(_00657_),
    .X(_10151_));
 sky130_fd_sc_hd__mux4_2 _24283_ (.A0(\w[35][18] ),
    .A1(\w[33][18] ),
    .A2(\w[39][18] ),
    .A3(\w[37][18] ),
    .S0(net361),
    .S1(net311),
    .X(_10152_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_522 ();
 sky130_fd_sc_hd__mux4_2 _24285_ (.A0(\w[43][18] ),
    .A1(\w[41][18] ),
    .A2(\w[47][18] ),
    .A3(\w[45][18] ),
    .S0(net363),
    .S1(net311),
    .X(_10154_));
 sky130_fd_sc_hd__mux4_2 _24286_ (.A0(_10150_),
    .A1(_10151_),
    .A2(_10152_),
    .A3(_10154_),
    .S0(net334),
    .S1(net327),
    .X(_10155_));
 sky130_fd_sc_hd__mux2i_1 _24287_ (.A0(_10149_),
    .A1(_10155_),
    .S(net293),
    .Y(_10156_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_521 ();
 sky130_fd_sc_hd__nand2_1 _24289_ (.A(net347),
    .B(\w[1][18] ),
    .Y(_10158_));
 sky130_fd_sc_hd__o21ai_0 _24290_ (.A1(net285),
    .A2(_10156_),
    .B1(_10158_),
    .Y(_00041_));
 sky130_fd_sc_hd__mux4_2 _24291_ (.A0(\w[19][19] ),
    .A1(\w[17][19] ),
    .A2(\w[23][19] ),
    .A3(\w[21][19] ),
    .S0(net361),
    .S1(net311),
    .X(_10159_));
 sky130_fd_sc_hd__mux4_2 _24292_ (.A0(\w[27][19] ),
    .A1(\w[25][19] ),
    .A2(\w[31][19] ),
    .A3(\w[29][19] ),
    .S0(net361),
    .S1(net311),
    .X(_10160_));
 sky130_fd_sc_hd__mux4_2 _24293_ (.A0(\w[3][19] ),
    .A1(\w[1][19] ),
    .A2(\w[7][19] ),
    .A3(\w[5][19] ),
    .S0(net361),
    .S1(net311),
    .X(_10161_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_520 ();
 sky130_fd_sc_hd__mux4_2 _24295_ (.A0(\w[11][19] ),
    .A1(\w[9][19] ),
    .A2(\w[15][19] ),
    .A3(\w[13][19] ),
    .S0(net361),
    .S1(net311),
    .X(_10163_));
 sky130_fd_sc_hd__mux4_2 _24296_ (.A0(_10159_),
    .A1(_10160_),
    .A2(_10161_),
    .A3(_10163_),
    .S0(net337),
    .S1(net329),
    .X(_10164_));
 sky130_fd_sc_hd__mux4_2 _24297_ (.A0(\w[51][19] ),
    .A1(\w[49][19] ),
    .A2(\w[55][19] ),
    .A3(\w[53][19] ),
    .S0(net363),
    .S1(_00657_),
    .X(_10165_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_519 ();
 sky130_fd_sc_hd__mux4_2 _24299_ (.A0(\w[59][19] ),
    .A1(\w[57][19] ),
    .A2(\w[63][19] ),
    .A3(\w[61][19] ),
    .S0(net363),
    .S1(_00657_),
    .X(_10167_));
 sky130_fd_sc_hd__mux4_2 _24300_ (.A0(\w[35][19] ),
    .A1(\w[33][19] ),
    .A2(\w[39][19] ),
    .A3(\w[37][19] ),
    .S0(net363),
    .S1(_00657_),
    .X(_10168_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_518 ();
 sky130_fd_sc_hd__mux4_2 _24302_ (.A0(\w[43][19] ),
    .A1(\w[41][19] ),
    .A2(\w[47][19] ),
    .A3(\w[45][19] ),
    .S0(net363),
    .S1(_00657_),
    .X(_10170_));
 sky130_fd_sc_hd__mux4_2 _24303_ (.A0(_10165_),
    .A1(_10167_),
    .A2(_10168_),
    .A3(_10170_),
    .S0(net338),
    .S1(_09857_),
    .X(_10171_));
 sky130_fd_sc_hd__mux2i_1 _24304_ (.A0(_10164_),
    .A1(_10171_),
    .S(net293),
    .Y(_10172_));
 sky130_fd_sc_hd__nand2_1 _24305_ (.A(net347),
    .B(\w[1][19] ),
    .Y(_10173_));
 sky130_fd_sc_hd__o21ai_0 _24306_ (.A1(net285),
    .A2(_10172_),
    .B1(_10173_),
    .Y(_00042_));
 sky130_fd_sc_hd__mux4_2 _24307_ (.A0(\w[19][20] ),
    .A1(\w[17][20] ),
    .A2(\w[23][20] ),
    .A3(\w[21][20] ),
    .S0(net361),
    .S1(net311),
    .X(_10174_));
 sky130_fd_sc_hd__mux4_2 _24308_ (.A0(\w[27][20] ),
    .A1(\w[25][20] ),
    .A2(\w[31][20] ),
    .A3(\w[29][20] ),
    .S0(net361),
    .S1(net311),
    .X(_10175_));
 sky130_fd_sc_hd__mux4_2 _24309_ (.A0(\w[3][20] ),
    .A1(\w[1][20] ),
    .A2(\w[7][20] ),
    .A3(\w[5][20] ),
    .S0(net361),
    .S1(net311),
    .X(_10176_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_517 ();
 sky130_fd_sc_hd__mux4_2 _24311_ (.A0(\w[11][20] ),
    .A1(\w[9][20] ),
    .A2(\w[15][20] ),
    .A3(\w[13][20] ),
    .S0(net361),
    .S1(net311),
    .X(_10178_));
 sky130_fd_sc_hd__mux4_2 _24312_ (.A0(_10174_),
    .A1(_10175_),
    .A2(_10176_),
    .A3(_10178_),
    .S0(net337),
    .S1(net329),
    .X(_10179_));
 sky130_fd_sc_hd__mux4_2 _24313_ (.A0(\w[51][20] ),
    .A1(\w[49][20] ),
    .A2(\w[55][20] ),
    .A3(\w[53][20] ),
    .S0(net364),
    .S1(net312),
    .X(_10180_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_516 ();
 sky130_fd_sc_hd__mux4_2 _24315_ (.A0(\w[59][20] ),
    .A1(\w[57][20] ),
    .A2(\w[63][20] ),
    .A3(\w[61][20] ),
    .S0(net364),
    .S1(net312),
    .X(_10182_));
 sky130_fd_sc_hd__mux4_2 _24316_ (.A0(\w[35][20] ),
    .A1(\w[33][20] ),
    .A2(\w[39][20] ),
    .A3(\w[37][20] ),
    .S0(net364),
    .S1(net312),
    .X(_10183_));
 sky130_fd_sc_hd__mux4_2 _24317_ (.A0(\w[43][20] ),
    .A1(\w[41][20] ),
    .A2(\w[47][20] ),
    .A3(\w[45][20] ),
    .S0(net364),
    .S1(net312),
    .X(_10184_));
 sky130_fd_sc_hd__mux4_2 _24318_ (.A0(_10180_),
    .A1(_10182_),
    .A2(_10183_),
    .A3(_10184_),
    .S0(_09854_),
    .S1(net331),
    .X(_10185_));
 sky130_fd_sc_hd__mux2i_1 _24319_ (.A0(_10179_),
    .A1(_10185_),
    .S(net293),
    .Y(_10186_));
 sky130_fd_sc_hd__nand2_1 _24320_ (.A(net347),
    .B(\w[1][20] ),
    .Y(_10187_));
 sky130_fd_sc_hd__o21ai_2 _24321_ (.A1(net285),
    .A2(_10186_),
    .B1(_10187_),
    .Y(_00044_));
 sky130_fd_sc_hd__mux4_2 _24322_ (.A0(\w[19][21] ),
    .A1(\w[17][21] ),
    .A2(\w[23][21] ),
    .A3(\w[21][21] ),
    .S0(net361),
    .S1(net311),
    .X(_10188_));
 sky130_fd_sc_hd__mux4_2 _24323_ (.A0(\w[27][21] ),
    .A1(\w[25][21] ),
    .A2(\w[31][21] ),
    .A3(\w[29][21] ),
    .S0(net361),
    .S1(net311),
    .X(_10189_));
 sky130_fd_sc_hd__mux4_2 _24324_ (.A0(\w[3][21] ),
    .A1(\w[1][21] ),
    .A2(\w[7][21] ),
    .A3(\w[5][21] ),
    .S0(net361),
    .S1(net311),
    .X(_10190_));
 sky130_fd_sc_hd__mux4_2 _24325_ (.A0(\w[11][21] ),
    .A1(\w[9][21] ),
    .A2(\w[15][21] ),
    .A3(\w[13][21] ),
    .S0(net361),
    .S1(net311),
    .X(_10191_));
 sky130_fd_sc_hd__mux4_2 _24326_ (.A0(_10188_),
    .A1(_10189_),
    .A2(_10190_),
    .A3(_10191_),
    .S0(net337),
    .S1(net329),
    .X(_10192_));
 sky130_fd_sc_hd__mux4_2 _24327_ (.A0(\w[51][21] ),
    .A1(\w[49][21] ),
    .A2(\w[55][21] ),
    .A3(\w[53][21] ),
    .S0(net363),
    .S1(net311),
    .X(_10193_));
 sky130_fd_sc_hd__mux4_2 _24328_ (.A0(\w[59][21] ),
    .A1(\w[57][21] ),
    .A2(\w[63][21] ),
    .A3(\w[61][21] ),
    .S0(net363),
    .S1(net311),
    .X(_10194_));
 sky130_fd_sc_hd__mux4_2 _24329_ (.A0(\w[35][21] ),
    .A1(\w[33][21] ),
    .A2(\w[39][21] ),
    .A3(\w[37][21] ),
    .S0(net363),
    .S1(net311),
    .X(_10195_));
 sky130_fd_sc_hd__mux4_2 _24330_ (.A0(\w[43][21] ),
    .A1(\w[41][21] ),
    .A2(\w[47][21] ),
    .A3(\w[45][21] ),
    .S0(net363),
    .S1(net311),
    .X(_10196_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_515 ();
 sky130_fd_sc_hd__mux4_2 _24332_ (.A0(_10193_),
    .A1(_10194_),
    .A2(_10195_),
    .A3(_10196_),
    .S0(net334),
    .S1(net327),
    .X(_10198_));
 sky130_fd_sc_hd__mux2i_1 _24333_ (.A0(_10192_),
    .A1(_10198_),
    .S(net293),
    .Y(_10199_));
 sky130_fd_sc_hd__nand2_1 _24334_ (.A(net347),
    .B(\w[1][21] ),
    .Y(_10200_));
 sky130_fd_sc_hd__o21ai_1 _24335_ (.A1(net285),
    .A2(_10199_),
    .B1(_10200_),
    .Y(_00045_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_514 ();
 sky130_fd_sc_hd__mux4_2 _24337_ (.A0(\w[19][22] ),
    .A1(\w[17][22] ),
    .A2(\w[23][22] ),
    .A3(\w[21][22] ),
    .S0(net361),
    .S1(net311),
    .X(_10202_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_513 ();
 sky130_fd_sc_hd__mux4_2 _24339_ (.A0(\w[27][22] ),
    .A1(\w[25][22] ),
    .A2(\w[31][22] ),
    .A3(\w[29][22] ),
    .S0(net361),
    .S1(net311),
    .X(_10204_));
 sky130_fd_sc_hd__mux4_2 _24340_ (.A0(\w[3][22] ),
    .A1(\w[1][22] ),
    .A2(\w[7][22] ),
    .A3(\w[5][22] ),
    .S0(net361),
    .S1(net311),
    .X(_10205_));
 sky130_fd_sc_hd__mux4_2 _24341_ (.A0(\w[11][22] ),
    .A1(\w[9][22] ),
    .A2(\w[15][22] ),
    .A3(\w[13][22] ),
    .S0(net361),
    .S1(net311),
    .X(_10206_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_512 ();
 sky130_fd_sc_hd__mux4_2 _24343_ (.A0(_10202_),
    .A1(_10204_),
    .A2(_10205_),
    .A3(_10206_),
    .S0(net337),
    .S1(net329),
    .X(_10208_));
 sky130_fd_sc_hd__mux4_2 _24344_ (.A0(\w[51][22] ),
    .A1(\w[49][22] ),
    .A2(\w[55][22] ),
    .A3(\w[53][22] ),
    .S0(net363),
    .S1(net311),
    .X(_10209_));
 sky130_fd_sc_hd__mux4_2 _24345_ (.A0(\w[59][22] ),
    .A1(\w[57][22] ),
    .A2(\w[63][22] ),
    .A3(\w[61][22] ),
    .S0(net363),
    .S1(net311),
    .X(_10210_));
 sky130_fd_sc_hd__mux4_2 _24346_ (.A0(\w[35][22] ),
    .A1(\w[33][22] ),
    .A2(\w[39][22] ),
    .A3(\w[37][22] ),
    .S0(net363),
    .S1(net311),
    .X(_10211_));
 sky130_fd_sc_hd__mux4_2 _24347_ (.A0(\w[43][22] ),
    .A1(\w[41][22] ),
    .A2(\w[47][22] ),
    .A3(\w[45][22] ),
    .S0(net363),
    .S1(net311),
    .X(_10212_));
 sky130_fd_sc_hd__mux4_2 _24348_ (.A0(_10209_),
    .A1(_10210_),
    .A2(_10211_),
    .A3(_10212_),
    .S0(net334),
    .S1(net327),
    .X(_10213_));
 sky130_fd_sc_hd__mux2i_1 _24349_ (.A0(_10208_),
    .A1(_10213_),
    .S(net293),
    .Y(_10214_));
 sky130_fd_sc_hd__nand2_1 _24350_ (.A(net347),
    .B(\w[1][22] ),
    .Y(_10215_));
 sky130_fd_sc_hd__o21ai_1 _24351_ (.A1(net285),
    .A2(_10214_),
    .B1(_10215_),
    .Y(_00046_));
 sky130_fd_sc_hd__mux4_2 _24352_ (.A0(\w[19][23] ),
    .A1(\w[17][23] ),
    .A2(\w[23][23] ),
    .A3(\w[21][23] ),
    .S0(net357),
    .S1(net308),
    .X(_10216_));
 sky130_fd_sc_hd__mux4_2 _24353_ (.A0(\w[27][23] ),
    .A1(\w[25][23] ),
    .A2(\w[31][23] ),
    .A3(\w[29][23] ),
    .S0(net357),
    .S1(net308),
    .X(_10217_));
 sky130_fd_sc_hd__mux4_2 _24354_ (.A0(\w[3][23] ),
    .A1(\w[1][23] ),
    .A2(\w[7][23] ),
    .A3(\w[5][23] ),
    .S0(net357),
    .S1(net308),
    .X(_10218_));
 sky130_fd_sc_hd__mux4_2 _24355_ (.A0(\w[11][23] ),
    .A1(\w[9][23] ),
    .A2(\w[15][23] ),
    .A3(\w[13][23] ),
    .S0(net357),
    .S1(net308),
    .X(_10219_));
 sky130_fd_sc_hd__mux4_2 _24356_ (.A0(_10216_),
    .A1(_10217_),
    .A2(_10218_),
    .A3(_10219_),
    .S0(net332),
    .S1(net331),
    .X(_10220_));
 sky130_fd_sc_hd__mux4_2 _24357_ (.A0(\w[51][23] ),
    .A1(\w[49][23] ),
    .A2(\w[55][23] ),
    .A3(\w[53][23] ),
    .S0(net360),
    .S1(net308),
    .X(_10221_));
 sky130_fd_sc_hd__mux4_2 _24358_ (.A0(\w[59][23] ),
    .A1(\w[57][23] ),
    .A2(\w[63][23] ),
    .A3(\w[61][23] ),
    .S0(net360),
    .S1(net308),
    .X(_10222_));
 sky130_fd_sc_hd__mux4_2 _24359_ (.A0(\w[35][23] ),
    .A1(\w[33][23] ),
    .A2(\w[39][23] ),
    .A3(\w[37][23] ),
    .S0(net360),
    .S1(net308),
    .X(_10223_));
 sky130_fd_sc_hd__mux4_2 _24360_ (.A0(\w[43][23] ),
    .A1(\w[41][23] ),
    .A2(\w[47][23] ),
    .A3(\w[45][23] ),
    .S0(net360),
    .S1(net308),
    .X(_10224_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_511 ();
 sky130_fd_sc_hd__mux4_2 _24362_ (.A0(_10221_),
    .A1(_10222_),
    .A2(_10223_),
    .A3(_10224_),
    .S0(net335),
    .S1(net330),
    .X(_10226_));
 sky130_fd_sc_hd__mux2i_1 _24363_ (.A0(_10220_),
    .A1(_10226_),
    .S(net295),
    .Y(_10227_));
 sky130_fd_sc_hd__nand2_2 _24364_ (.A(net349),
    .B(\w[1][23] ),
    .Y(_10228_));
 sky130_fd_sc_hd__o21ai_4 _24365_ (.A1(net287),
    .A2(_10227_),
    .B1(_10228_),
    .Y(_00047_));
 sky130_fd_sc_hd__mux4_2 _24366_ (.A0(\w[19][24] ),
    .A1(\w[17][24] ),
    .A2(\w[23][24] ),
    .A3(\w[21][24] ),
    .S0(net359),
    .S1(net309),
    .X(_10229_));
 sky130_fd_sc_hd__mux4_2 _24367_ (.A0(\w[27][24] ),
    .A1(\w[25][24] ),
    .A2(\w[31][24] ),
    .A3(\w[29][24] ),
    .S0(net359),
    .S1(net309),
    .X(_10230_));
 sky130_fd_sc_hd__mux4_2 _24368_ (.A0(\w[3][24] ),
    .A1(\w[1][24] ),
    .A2(\w[7][24] ),
    .A3(\w[5][24] ),
    .S0(net359),
    .S1(net309),
    .X(_10231_));
 sky130_fd_sc_hd__mux4_2 _24369_ (.A0(\w[11][24] ),
    .A1(\w[9][24] ),
    .A2(\w[15][24] ),
    .A3(\w[13][24] ),
    .S0(net359),
    .S1(net309),
    .X(_10232_));
 sky130_fd_sc_hd__mux4_2 _24370_ (.A0(_10229_),
    .A1(_10230_),
    .A2(_10231_),
    .A3(_10232_),
    .S0(net333),
    .S1(net327),
    .X(_10233_));
 sky130_fd_sc_hd__mux4_2 _24371_ (.A0(\w[51][24] ),
    .A1(\w[49][24] ),
    .A2(\w[55][24] ),
    .A3(\w[53][24] ),
    .S0(net360),
    .S1(net308),
    .X(_10234_));
 sky130_fd_sc_hd__mux4_2 _24372_ (.A0(\w[59][24] ),
    .A1(\w[57][24] ),
    .A2(\w[63][24] ),
    .A3(\w[61][24] ),
    .S0(net360),
    .S1(net308),
    .X(_10235_));
 sky130_fd_sc_hd__mux4_2 _24373_ (.A0(\w[35][24] ),
    .A1(\w[33][24] ),
    .A2(\w[39][24] ),
    .A3(\w[37][24] ),
    .S0(net360),
    .S1(net308),
    .X(_10236_));
 sky130_fd_sc_hd__mux4_2 _24374_ (.A0(\w[43][24] ),
    .A1(\w[41][24] ),
    .A2(\w[47][24] ),
    .A3(\w[45][24] ),
    .S0(net360),
    .S1(net308),
    .X(_10237_));
 sky130_fd_sc_hd__mux4_2 _24375_ (.A0(_10234_),
    .A1(_10235_),
    .A2(_10236_),
    .A3(_10237_),
    .S0(net335),
    .S1(net328),
    .X(_10238_));
 sky130_fd_sc_hd__mux2i_1 _24376_ (.A0(_10233_),
    .A1(_10238_),
    .S(net292),
    .Y(_10239_));
 sky130_fd_sc_hd__nand2_2 _24377_ (.A(net347),
    .B(\w[1][24] ),
    .Y(_10240_));
 sky130_fd_sc_hd__o21ai_4 _24378_ (.A1(net285),
    .A2(_10239_),
    .B1(_10240_),
    .Y(_00048_));
 sky130_fd_sc_hd__mux4_2 _24379_ (.A0(\w[19][25] ),
    .A1(\w[17][25] ),
    .A2(\w[23][25] ),
    .A3(\w[21][25] ),
    .S0(net363),
    .S1(net311),
    .X(_10241_));
 sky130_fd_sc_hd__mux4_2 _24380_ (.A0(\w[27][25] ),
    .A1(\w[25][25] ),
    .A2(\w[31][25] ),
    .A3(\w[29][25] ),
    .S0(net363),
    .S1(net311),
    .X(_10242_));
 sky130_fd_sc_hd__mux4_2 _24381_ (.A0(\w[3][25] ),
    .A1(\w[1][25] ),
    .A2(\w[7][25] ),
    .A3(\w[5][25] ),
    .S0(net363),
    .S1(net311),
    .X(_10243_));
 sky130_fd_sc_hd__mux4_2 _24382_ (.A0(\w[11][25] ),
    .A1(\w[9][25] ),
    .A2(\w[15][25] ),
    .A3(\w[13][25] ),
    .S0(net363),
    .S1(net311),
    .X(_10244_));
 sky130_fd_sc_hd__mux4_2 _24383_ (.A0(_10241_),
    .A1(_10242_),
    .A2(_10243_),
    .A3(_10244_),
    .S0(net334),
    .S1(net327),
    .X(_10245_));
 sky130_fd_sc_hd__mux4_2 _24384_ (.A0(\w[51][25] ),
    .A1(\w[49][25] ),
    .A2(\w[55][25] ),
    .A3(\w[53][25] ),
    .S0(net359),
    .S1(net309),
    .X(_10246_));
 sky130_fd_sc_hd__mux4_2 _24385_ (.A0(\w[59][25] ),
    .A1(\w[57][25] ),
    .A2(\w[63][25] ),
    .A3(\w[61][25] ),
    .S0(net359),
    .S1(net309),
    .X(_10247_));
 sky130_fd_sc_hd__mux4_2 _24386_ (.A0(\w[35][25] ),
    .A1(\w[33][25] ),
    .A2(\w[39][25] ),
    .A3(\w[37][25] ),
    .S0(net359),
    .S1(net309),
    .X(_10248_));
 sky130_fd_sc_hd__mux4_2 _24387_ (.A0(\w[43][25] ),
    .A1(\w[41][25] ),
    .A2(\w[47][25] ),
    .A3(\w[45][25] ),
    .S0(net359),
    .S1(net309),
    .X(_10249_));
 sky130_fd_sc_hd__mux4_2 _24388_ (.A0(_10246_),
    .A1(_10247_),
    .A2(_10248_),
    .A3(_10249_),
    .S0(net333),
    .S1(net327),
    .X(_10250_));
 sky130_fd_sc_hd__mux2i_1 _24389_ (.A0(_10245_),
    .A1(_10250_),
    .S(net292),
    .Y(_10251_));
 sky130_fd_sc_hd__nand2_1 _24390_ (.A(net347),
    .B(\w[1][25] ),
    .Y(_10252_));
 sky130_fd_sc_hd__o21ai_2 _24391_ (.A1(net285),
    .A2(_10251_),
    .B1(_10252_),
    .Y(_00049_));
 sky130_fd_sc_hd__mux4_2 _24392_ (.A0(\w[19][26] ),
    .A1(\w[17][26] ),
    .A2(\w[23][26] ),
    .A3(\w[21][26] ),
    .S0(net357),
    .S1(net312),
    .X(_10253_));
 sky130_fd_sc_hd__mux4_2 _24393_ (.A0(\w[27][26] ),
    .A1(\w[25][26] ),
    .A2(\w[31][26] ),
    .A3(\w[29][26] ),
    .S0(net357),
    .S1(net312),
    .X(_10254_));
 sky130_fd_sc_hd__mux4_2 _24394_ (.A0(\w[3][26] ),
    .A1(\w[1][26] ),
    .A2(\w[7][26] ),
    .A3(\w[5][26] ),
    .S0(net357),
    .S1(net312),
    .X(_10255_));
 sky130_fd_sc_hd__mux4_2 _24395_ (.A0(\w[11][26] ),
    .A1(\w[9][26] ),
    .A2(\w[15][26] ),
    .A3(\w[13][26] ),
    .S0(net357),
    .S1(net312),
    .X(_10256_));
 sky130_fd_sc_hd__mux4_2 _24396_ (.A0(_10253_),
    .A1(_10254_),
    .A2(_10255_),
    .A3(_10256_),
    .S0(net332),
    .S1(net331),
    .X(_10257_));
 sky130_fd_sc_hd__mux4_2 _24397_ (.A0(\w[51][26] ),
    .A1(\w[49][26] ),
    .A2(\w[55][26] ),
    .A3(\w[53][26] ),
    .S0(net364),
    .S1(net312),
    .X(_10258_));
 sky130_fd_sc_hd__mux4_2 _24398_ (.A0(\w[59][26] ),
    .A1(\w[57][26] ),
    .A2(\w[63][26] ),
    .A3(\w[61][26] ),
    .S0(net364),
    .S1(net312),
    .X(_10259_));
 sky130_fd_sc_hd__mux4_2 _24399_ (.A0(\w[35][26] ),
    .A1(\w[33][26] ),
    .A2(\w[39][26] ),
    .A3(\w[37][26] ),
    .S0(net364),
    .S1(net312),
    .X(_10260_));
 sky130_fd_sc_hd__mux4_2 _24400_ (.A0(\w[43][26] ),
    .A1(\w[41][26] ),
    .A2(\w[47][26] ),
    .A3(\w[45][26] ),
    .S0(net364),
    .S1(net312),
    .X(_10261_));
 sky130_fd_sc_hd__mux4_2 _24401_ (.A0(_10258_),
    .A1(_10259_),
    .A2(_10260_),
    .A3(_10261_),
    .S0(net332),
    .S1(net330),
    .X(_10262_));
 sky130_fd_sc_hd__mux2i_1 _24402_ (.A0(_10257_),
    .A1(_10262_),
    .S(net295),
    .Y(_10263_));
 sky130_fd_sc_hd__nand2_2 _24403_ (.A(net349),
    .B(\w[1][26] ),
    .Y(_10264_));
 sky130_fd_sc_hd__o21ai_4 _24404_ (.A1(net287),
    .A2(_10263_),
    .B1(_10264_),
    .Y(_00050_));
 sky130_fd_sc_hd__mux4_2 _24405_ (.A0(\w[19][27] ),
    .A1(\w[17][27] ),
    .A2(\w[23][27] ),
    .A3(\w[21][27] ),
    .S0(net358),
    .S1(net310),
    .X(_10265_));
 sky130_fd_sc_hd__mux4_2 _24406_ (.A0(\w[27][27] ),
    .A1(\w[25][27] ),
    .A2(\w[31][27] ),
    .A3(\w[29][27] ),
    .S0(net358),
    .S1(net310),
    .X(_10266_));
 sky130_fd_sc_hd__mux4_2 _24407_ (.A0(\w[3][27] ),
    .A1(\w[1][27] ),
    .A2(\w[7][27] ),
    .A3(\w[5][27] ),
    .S0(net358),
    .S1(net310),
    .X(_10267_));
 sky130_fd_sc_hd__mux4_2 _24408_ (.A0(\w[11][27] ),
    .A1(\w[9][27] ),
    .A2(\w[15][27] ),
    .A3(\w[13][27] ),
    .S0(net358),
    .S1(net310),
    .X(_10268_));
 sky130_fd_sc_hd__mux4_2 _24409_ (.A0(_10265_),
    .A1(_10266_),
    .A2(_10267_),
    .A3(_10268_),
    .S0(net336),
    .S1(net326),
    .X(_10269_));
 sky130_fd_sc_hd__mux4_2 _24410_ (.A0(\w[51][27] ),
    .A1(\w[49][27] ),
    .A2(\w[55][27] ),
    .A3(\w[53][27] ),
    .S0(net360),
    .S1(net308),
    .X(_10270_));
 sky130_fd_sc_hd__mux4_2 _24411_ (.A0(\w[59][27] ),
    .A1(\w[57][27] ),
    .A2(\w[63][27] ),
    .A3(\w[61][27] ),
    .S0(net360),
    .S1(net308),
    .X(_10271_));
 sky130_fd_sc_hd__mux4_2 _24412_ (.A0(\w[35][27] ),
    .A1(\w[33][27] ),
    .A2(\w[39][27] ),
    .A3(\w[37][27] ),
    .S0(net360),
    .S1(net308),
    .X(_10272_));
 sky130_fd_sc_hd__mux4_2 _24413_ (.A0(\w[43][27] ),
    .A1(\w[41][27] ),
    .A2(\w[47][27] ),
    .A3(\w[45][27] ),
    .S0(net360),
    .S1(net308),
    .X(_10273_));
 sky130_fd_sc_hd__mux4_2 _24414_ (.A0(_10270_),
    .A1(_10271_),
    .A2(_10272_),
    .A3(_10273_),
    .S0(net335),
    .S1(net328),
    .X(_10274_));
 sky130_fd_sc_hd__mux2i_1 _24415_ (.A0(_10269_),
    .A1(_10274_),
    .S(net292),
    .Y(_10275_));
 sky130_fd_sc_hd__nand2_2 _24416_ (.A(net347),
    .B(\w[1][27] ),
    .Y(_10276_));
 sky130_fd_sc_hd__o21ai_4 _24417_ (.A1(net285),
    .A2(_10275_),
    .B1(_10276_),
    .Y(_00051_));
 sky130_fd_sc_hd__mux4_2 _24418_ (.A0(\w[19][28] ),
    .A1(\w[17][28] ),
    .A2(\w[23][28] ),
    .A3(\w[21][28] ),
    .S0(net357),
    .S1(net308),
    .X(_10277_));
 sky130_fd_sc_hd__mux4_2 _24419_ (.A0(\w[27][28] ),
    .A1(\w[25][28] ),
    .A2(\w[31][28] ),
    .A3(\w[29][28] ),
    .S0(net357),
    .S1(net308),
    .X(_10278_));
 sky130_fd_sc_hd__mux4_2 _24420_ (.A0(\w[3][28] ),
    .A1(\w[1][28] ),
    .A2(\w[7][28] ),
    .A3(\w[5][28] ),
    .S0(net357),
    .S1(net308),
    .X(_10279_));
 sky130_fd_sc_hd__mux4_2 _24421_ (.A0(\w[11][28] ),
    .A1(\w[9][28] ),
    .A2(\w[15][28] ),
    .A3(\w[13][28] ),
    .S0(net357),
    .S1(net308),
    .X(_10280_));
 sky130_fd_sc_hd__mux4_2 _24422_ (.A0(_10277_),
    .A1(_10278_),
    .A2(_10279_),
    .A3(_10280_),
    .S0(net332),
    .S1(net331),
    .X(_10281_));
 sky130_fd_sc_hd__mux4_2 _24423_ (.A0(\w[51][28] ),
    .A1(\w[49][28] ),
    .A2(\w[55][28] ),
    .A3(\w[53][28] ),
    .S0(net364),
    .S1(net308),
    .X(_10282_));
 sky130_fd_sc_hd__mux4_2 _24424_ (.A0(\w[59][28] ),
    .A1(\w[57][28] ),
    .A2(\w[63][28] ),
    .A3(\w[61][28] ),
    .S0(net364),
    .S1(net308),
    .X(_10283_));
 sky130_fd_sc_hd__mux4_2 _24425_ (.A0(\w[35][28] ),
    .A1(\w[33][28] ),
    .A2(\w[39][28] ),
    .A3(\w[37][28] ),
    .S0(net364),
    .S1(net308),
    .X(_10284_));
 sky130_fd_sc_hd__mux4_2 _24426_ (.A0(\w[43][28] ),
    .A1(\w[41][28] ),
    .A2(\w[47][28] ),
    .A3(\w[45][28] ),
    .S0(net364),
    .S1(net308),
    .X(_10285_));
 sky130_fd_sc_hd__mux4_2 _24427_ (.A0(_10282_),
    .A1(_10283_),
    .A2(_10284_),
    .A3(_10285_),
    .S0(net332),
    .S1(net330),
    .X(_10286_));
 sky130_fd_sc_hd__mux2i_2 _24428_ (.A0(_10281_),
    .A1(_10286_),
    .S(net295),
    .Y(_10287_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_510 ();
 sky130_fd_sc_hd__nand2_2 _24430_ (.A(net349),
    .B(\w[1][28] ),
    .Y(_10289_));
 sky130_fd_sc_hd__o21ai_4 _24431_ (.A1(net287),
    .A2(_10287_),
    .B1(_10289_),
    .Y(_00052_));
 sky130_fd_sc_hd__mux4_2 _24432_ (.A0(\w[19][29] ),
    .A1(\w[17][29] ),
    .A2(\w[23][29] ),
    .A3(\w[21][29] ),
    .S0(net357),
    .S1(net312),
    .X(_10290_));
 sky130_fd_sc_hd__mux4_2 _24433_ (.A0(\w[27][29] ),
    .A1(\w[25][29] ),
    .A2(\w[31][29] ),
    .A3(\w[29][29] ),
    .S0(net357),
    .S1(net312),
    .X(_10291_));
 sky130_fd_sc_hd__mux4_2 _24434_ (.A0(\w[3][29] ),
    .A1(\w[1][29] ),
    .A2(\w[7][29] ),
    .A3(\w[5][29] ),
    .S0(net357),
    .S1(net312),
    .X(_10292_));
 sky130_fd_sc_hd__mux4_2 _24435_ (.A0(\w[11][29] ),
    .A1(\w[9][29] ),
    .A2(\w[15][29] ),
    .A3(\w[13][29] ),
    .S0(net357),
    .S1(net312),
    .X(_10293_));
 sky130_fd_sc_hd__mux4_2 _24436_ (.A0(_10290_),
    .A1(_10291_),
    .A2(_10292_),
    .A3(_10293_),
    .S0(net332),
    .S1(net331),
    .X(_10294_));
 sky130_fd_sc_hd__mux4_2 _24437_ (.A0(\w[51][29] ),
    .A1(\w[49][29] ),
    .A2(\w[55][29] ),
    .A3(\w[53][29] ),
    .S0(net364),
    .S1(net308),
    .X(_10295_));
 sky130_fd_sc_hd__mux4_2 _24438_ (.A0(\w[59][29] ),
    .A1(\w[57][29] ),
    .A2(\w[63][29] ),
    .A3(\w[61][29] ),
    .S0(net364),
    .S1(net308),
    .X(_10296_));
 sky130_fd_sc_hd__mux4_2 _24439_ (.A0(\w[35][29] ),
    .A1(\w[33][29] ),
    .A2(\w[39][29] ),
    .A3(\w[37][29] ),
    .S0(net364),
    .S1(net308),
    .X(_10297_));
 sky130_fd_sc_hd__mux4_2 _24440_ (.A0(\w[43][29] ),
    .A1(\w[41][29] ),
    .A2(\w[47][29] ),
    .A3(\w[45][29] ),
    .S0(net364),
    .S1(net308),
    .X(_10298_));
 sky130_fd_sc_hd__mux4_2 _24441_ (.A0(_10295_),
    .A1(_10296_),
    .A2(_10297_),
    .A3(_10298_),
    .S0(net332),
    .S1(net330),
    .X(_10299_));
 sky130_fd_sc_hd__mux2i_1 _24442_ (.A0(_10294_),
    .A1(_10299_),
    .S(net295),
    .Y(_10300_));
 sky130_fd_sc_hd__nand2_2 _24443_ (.A(net349),
    .B(\w[1][29] ),
    .Y(_10301_));
 sky130_fd_sc_hd__o21ai_4 _24444_ (.A1(net287),
    .A2(_10300_),
    .B1(_10301_),
    .Y(_00053_));
 sky130_fd_sc_hd__mux4_2 _24445_ (.A0(\w[19][30] ),
    .A1(\w[17][30] ),
    .A2(\w[23][30] ),
    .A3(\w[21][30] ),
    .S0(net357),
    .S1(net312),
    .X(_10302_));
 sky130_fd_sc_hd__mux4_2 _24446_ (.A0(\w[27][30] ),
    .A1(\w[25][30] ),
    .A2(\w[31][30] ),
    .A3(\w[29][30] ),
    .S0(net357),
    .S1(net312),
    .X(_10303_));
 sky130_fd_sc_hd__mux4_2 _24447_ (.A0(\w[3][30] ),
    .A1(\w[1][30] ),
    .A2(\w[7][30] ),
    .A3(\w[5][30] ),
    .S0(net357),
    .S1(net312),
    .X(_10304_));
 sky130_fd_sc_hd__mux4_2 _24448_ (.A0(\w[11][30] ),
    .A1(\w[9][30] ),
    .A2(\w[15][30] ),
    .A3(\w[13][30] ),
    .S0(net357),
    .S1(net312),
    .X(_10305_));
 sky130_fd_sc_hd__mux4_2 _24449_ (.A0(_10302_),
    .A1(_10303_),
    .A2(_10304_),
    .A3(_10305_),
    .S0(net332),
    .S1(net331),
    .X(_10306_));
 sky130_fd_sc_hd__mux4_2 _24450_ (.A0(\w[51][30] ),
    .A1(\w[49][30] ),
    .A2(\w[55][30] ),
    .A3(\w[53][30] ),
    .S0(net364),
    .S1(net312),
    .X(_10307_));
 sky130_fd_sc_hd__mux4_2 _24451_ (.A0(\w[59][30] ),
    .A1(\w[57][30] ),
    .A2(\w[63][30] ),
    .A3(\w[61][30] ),
    .S0(net364),
    .S1(net312),
    .X(_10308_));
 sky130_fd_sc_hd__mux4_2 _24452_ (.A0(\w[35][30] ),
    .A1(\w[33][30] ),
    .A2(\w[39][30] ),
    .A3(\w[37][30] ),
    .S0(net364),
    .S1(net312),
    .X(_10309_));
 sky130_fd_sc_hd__mux4_2 _24453_ (.A0(\w[43][30] ),
    .A1(\w[41][30] ),
    .A2(\w[47][30] ),
    .A3(\w[45][30] ),
    .S0(net364),
    .S1(net312),
    .X(_10310_));
 sky130_fd_sc_hd__mux4_2 _24454_ (.A0(_10307_),
    .A1(_10308_),
    .A2(_10309_),
    .A3(_10310_),
    .S0(net332),
    .S1(net331),
    .X(_10311_));
 sky130_fd_sc_hd__mux2i_1 _24455_ (.A0(_10306_),
    .A1(_10311_),
    .S(net295),
    .Y(_10312_));
 sky130_fd_sc_hd__nand2_2 _24456_ (.A(net349),
    .B(\w[1][30] ),
    .Y(_10313_));
 sky130_fd_sc_hd__o21ai_4 _24457_ (.A1(net287),
    .A2(_10312_),
    .B1(_10313_),
    .Y(_00055_));
 sky130_fd_sc_hd__mux4_2 _24458_ (.A0(\w[19][31] ),
    .A1(\w[17][31] ),
    .A2(\w[23][31] ),
    .A3(\w[21][31] ),
    .S0(net358),
    .S1(net310),
    .X(_10314_));
 sky130_fd_sc_hd__mux4_2 _24459_ (.A0(\w[27][31] ),
    .A1(\w[25][31] ),
    .A2(\w[31][31] ),
    .A3(\w[29][31] ),
    .S0(net358),
    .S1(net310),
    .X(_10315_));
 sky130_fd_sc_hd__mux4_2 _24460_ (.A0(\w[3][31] ),
    .A1(\w[1][31] ),
    .A2(\w[7][31] ),
    .A3(\w[5][31] ),
    .S0(net358),
    .S1(net310),
    .X(_10316_));
 sky130_fd_sc_hd__mux4_2 _24461_ (.A0(\w[11][31] ),
    .A1(\w[9][31] ),
    .A2(\w[15][31] ),
    .A3(\w[13][31] ),
    .S0(net358),
    .S1(net310),
    .X(_10317_));
 sky130_fd_sc_hd__mux4_2 _24462_ (.A0(_10314_),
    .A1(_10315_),
    .A2(_10316_),
    .A3(_10317_),
    .S0(net333),
    .S1(net326),
    .X(_10318_));
 sky130_fd_sc_hd__mux4_2 _24463_ (.A0(\w[51][31] ),
    .A1(\w[49][31] ),
    .A2(\w[55][31] ),
    .A3(\w[53][31] ),
    .S0(net358),
    .S1(net310),
    .X(_10319_));
 sky130_fd_sc_hd__mux4_2 _24464_ (.A0(\w[59][31] ),
    .A1(\w[57][31] ),
    .A2(\w[63][31] ),
    .A3(\w[61][31] ),
    .S0(net358),
    .S1(net310),
    .X(_10320_));
 sky130_fd_sc_hd__mux4_2 _24465_ (.A0(\w[35][31] ),
    .A1(\w[33][31] ),
    .A2(\w[39][31] ),
    .A3(\w[37][31] ),
    .S0(net358),
    .S1(net310),
    .X(_10321_));
 sky130_fd_sc_hd__mux4_2 _24466_ (.A0(\w[43][31] ),
    .A1(\w[41][31] ),
    .A2(\w[47][31] ),
    .A3(\w[45][31] ),
    .S0(net358),
    .S1(net310),
    .X(_10322_));
 sky130_fd_sc_hd__mux4_2 _24467_ (.A0(_10319_),
    .A1(_10320_),
    .A2(_10321_),
    .A3(_10322_),
    .S0(net336),
    .S1(net326),
    .X(_10323_));
 sky130_fd_sc_hd__mux2i_1 _24468_ (.A0(_10318_),
    .A1(_10323_),
    .S(net292),
    .Y(_10324_));
 sky130_fd_sc_hd__nand2_2 _24469_ (.A(net347),
    .B(\w[1][31] ),
    .Y(_10325_));
 sky130_fd_sc_hd__o21ai_4 _24470_ (.A1(net285),
    .A2(_10324_),
    .B1(_10325_),
    .Y(_00056_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_503 ();
 sky130_fd_sc_hd__mux4_2 _24478_ (.A0(\w[18][0] ),
    .A1(\w[16][0] ),
    .A2(\w[22][0] ),
    .A3(\w[20][0] ),
    .S0(net371),
    .S1(net307),
    .X(_10333_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_499 ();
 sky130_fd_sc_hd__mux4_2 _24483_ (.A0(\w[26][0] ),
    .A1(\w[24][0] ),
    .A2(\w[30][0] ),
    .A3(\w[28][0] ),
    .S0(net371),
    .S1(net307),
    .X(_10338_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_497 ();
 sky130_fd_sc_hd__mux4_2 _24486_ (.A0(\w[2][0] ),
    .A1(\w[0][0] ),
    .A2(\w[6][0] ),
    .A3(\w[4][0] ),
    .S0(net371),
    .S1(net307),
    .X(_10341_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_493 ();
 sky130_fd_sc_hd__mux4_2 _24491_ (.A0(\w[10][0] ),
    .A1(\w[8][0] ),
    .A2(\w[14][0] ),
    .A3(\w[12][0] ),
    .S0(net371),
    .S1(net307),
    .X(_10346_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_492 ();
 sky130_fd_sc_hd__xor2_4 _24493_ (.A(\count_hash1[3] ),
    .B(_12920_),
    .X(_10348_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_490 ();
 sky130_fd_sc_hd__nand3_4 _24496_ (.A(\count_hash1[3] ),
    .B(\count_hash1[2] ),
    .C(\count_hash1[1] ),
    .Y(_10351_));
 sky130_fd_sc_hd__xor2_4 _24497_ (.A(\count_hash1[4] ),
    .B(_10351_),
    .X(_10352_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_488 ();
 sky130_fd_sc_hd__mux4_2 _24500_ (.A0(_10333_),
    .A1(_10338_),
    .A2(_10341_),
    .A3(_10346_),
    .S0(net320),
    .S1(net316),
    .X(_10355_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_486 ();
 sky130_fd_sc_hd__mux4_2 _24503_ (.A0(\w[50][0] ),
    .A1(\w[48][0] ),
    .A2(\w[54][0] ),
    .A3(\w[52][0] ),
    .S0(net372),
    .S1(net303),
    .X(_10358_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_484 ();
 sky130_fd_sc_hd__mux4_2 _24506_ (.A0(\w[58][0] ),
    .A1(\w[56][0] ),
    .A2(\w[62][0] ),
    .A3(\w[60][0] ),
    .S0(net372),
    .S1(net303),
    .X(_10361_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_482 ();
 sky130_fd_sc_hd__mux4_2 _24509_ (.A0(\w[34][0] ),
    .A1(\w[32][0] ),
    .A2(\w[38][0] ),
    .A3(\w[36][0] ),
    .S0(net372),
    .S1(net303),
    .X(_10364_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_480 ();
 sky130_fd_sc_hd__mux4_2 _24512_ (.A0(\w[42][0] ),
    .A1(\w[40][0] ),
    .A2(\w[46][0] ),
    .A3(\w[44][0] ),
    .S0(net372),
    .S1(net303),
    .X(_10367_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_477 ();
 sky130_fd_sc_hd__mux4_2 _24516_ (.A0(_10358_),
    .A1(_10361_),
    .A2(_10364_),
    .A3(_10367_),
    .S0(net321),
    .S1(net317),
    .X(_10371_));
 sky130_fd_sc_hd__nand3_4 _24517_ (.A(\count_hash1[4] ),
    .B(\count_hash1[3] ),
    .C(_12920_),
    .Y(_10372_));
 sky130_fd_sc_hd__xnor2_4 _24518_ (.A(\count_hash1[5] ),
    .B(_10372_),
    .Y(_10373_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_474 ();
 sky130_fd_sc_hd__mux2i_1 _24522_ (.A0(_10355_),
    .A1(_10371_),
    .S(net290),
    .Y(_10377_));
 sky130_fd_sc_hd__nand2_1 _24523_ (.A(net348),
    .B(\w[0][0] ),
    .Y(_10378_));
 sky130_fd_sc_hd__o21ai_0 _24524_ (.A1(net287),
    .A2(_10377_),
    .B1(_10378_),
    .Y(_00000_));
 sky130_fd_sc_hd__mux4_2 _24525_ (.A0(\w[18][1] ),
    .A1(\w[16][1] ),
    .A2(\w[22][1] ),
    .A3(\w[20][1] ),
    .S0(net371),
    .S1(net307),
    .X(_10379_));
 sky130_fd_sc_hd__mux4_2 _24526_ (.A0(\w[26][1] ),
    .A1(\w[24][1] ),
    .A2(\w[30][1] ),
    .A3(\w[28][1] ),
    .S0(net372),
    .S1(net307),
    .X(_10380_));
 sky130_fd_sc_hd__mux4_2 _24527_ (.A0(\w[2][1] ),
    .A1(\w[0][1] ),
    .A2(\w[6][1] ),
    .A3(\w[4][1] ),
    .S0(net371),
    .S1(net307),
    .X(_10381_));
 sky130_fd_sc_hd__mux4_2 _24528_ (.A0(\w[10][1] ),
    .A1(\w[8][1] ),
    .A2(\w[14][1] ),
    .A3(\w[12][1] ),
    .S0(net371),
    .S1(net307),
    .X(_10382_));
 sky130_fd_sc_hd__mux4_2 _24529_ (.A0(_10379_),
    .A1(_10380_),
    .A2(_10381_),
    .A3(_10382_),
    .S0(net321),
    .S1(net317),
    .X(_10383_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_473 ();
 sky130_fd_sc_hd__mux4_2 _24531_ (.A0(\w[50][1] ),
    .A1(\w[48][1] ),
    .A2(\w[54][1] ),
    .A3(\w[52][1] ),
    .S0(net370),
    .S1(net306),
    .X(_10385_));
 sky130_fd_sc_hd__mux4_2 _24532_ (.A0(\w[58][1] ),
    .A1(\w[56][1] ),
    .A2(\w[62][1] ),
    .A3(\w[60][1] ),
    .S0(net370),
    .S1(net306),
    .X(_10386_));
 sky130_fd_sc_hd__mux4_2 _24533_ (.A0(\w[34][1] ),
    .A1(\w[32][1] ),
    .A2(\w[38][1] ),
    .A3(\w[36][1] ),
    .S0(net370),
    .S1(net306),
    .X(_10387_));
 sky130_fd_sc_hd__mux4_2 _24534_ (.A0(\w[42][1] ),
    .A1(\w[40][1] ),
    .A2(\w[46][1] ),
    .A3(\w[44][1] ),
    .S0(net370),
    .S1(net306),
    .X(_10388_));
 sky130_fd_sc_hd__mux4_2 _24535_ (.A0(_10385_),
    .A1(_10386_),
    .A2(_10387_),
    .A3(_10388_),
    .S0(net324),
    .S1(net315),
    .X(_10389_));
 sky130_fd_sc_hd__mux2i_1 _24536_ (.A0(_10383_),
    .A1(_10389_),
    .S(net289),
    .Y(_10390_));
 sky130_fd_sc_hd__nand2_1 _24537_ (.A(net348),
    .B(\w[0][1] ),
    .Y(_10391_));
 sky130_fd_sc_hd__o21ai_2 _24538_ (.A1(net286),
    .A2(_10390_),
    .B1(_10391_),
    .Y(_00011_));
 sky130_fd_sc_hd__mux4_2 _24539_ (.A0(\w[18][2] ),
    .A1(\w[16][2] ),
    .A2(\w[22][2] ),
    .A3(\w[20][2] ),
    .S0(net367),
    .S1(net303),
    .X(_10392_));
 sky130_fd_sc_hd__mux4_2 _24540_ (.A0(\w[26][2] ),
    .A1(\w[24][2] ),
    .A2(\w[30][2] ),
    .A3(\w[28][2] ),
    .S0(net367),
    .S1(net303),
    .X(_10393_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_472 ();
 sky130_fd_sc_hd__mux4_2 _24542_ (.A0(\w[2][2] ),
    .A1(\w[0][2] ),
    .A2(\w[6][2] ),
    .A3(\w[4][2] ),
    .S0(net367),
    .S1(net303),
    .X(_10395_));
 sky130_fd_sc_hd__mux4_2 _24543_ (.A0(\w[10][2] ),
    .A1(\w[8][2] ),
    .A2(\w[14][2] ),
    .A3(\w[12][2] ),
    .S0(net367),
    .S1(net303),
    .X(_10396_));
 sky130_fd_sc_hd__mux4_2 _24544_ (.A0(_10392_),
    .A1(_10393_),
    .A2(_10395_),
    .A3(_10396_),
    .S0(net322),
    .S1(net313),
    .X(_10397_));
 sky130_fd_sc_hd__mux4_2 _24545_ (.A0(\w[50][2] ),
    .A1(\w[48][2] ),
    .A2(\w[54][2] ),
    .A3(\w[52][2] ),
    .S0(net366),
    .S1(net306),
    .X(_10398_));
 sky130_fd_sc_hd__mux4_2 _24546_ (.A0(\w[58][2] ),
    .A1(\w[56][2] ),
    .A2(\w[62][2] ),
    .A3(\w[60][2] ),
    .S0(net366),
    .S1(net306),
    .X(_10399_));
 sky130_fd_sc_hd__mux4_2 _24547_ (.A0(\w[34][2] ),
    .A1(\w[32][2] ),
    .A2(\w[38][2] ),
    .A3(\w[36][2] ),
    .S0(net366),
    .S1(net306),
    .X(_10400_));
 sky130_fd_sc_hd__mux4_2 _24548_ (.A0(\w[42][2] ),
    .A1(\w[40][2] ),
    .A2(\w[46][2] ),
    .A3(\w[44][2] ),
    .S0(net366),
    .S1(net306),
    .X(_10401_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_471 ();
 sky130_fd_sc_hd__mux4_2 _24550_ (.A0(_10398_),
    .A1(_10399_),
    .A2(_10400_),
    .A3(_10401_),
    .S0(net323),
    .S1(net314),
    .X(_10403_));
 sky130_fd_sc_hd__mux2i_1 _24551_ (.A0(_10397_),
    .A1(_10403_),
    .S(net288),
    .Y(_10404_));
 sky130_fd_sc_hd__nand2_2 _24552_ (.A(net348),
    .B(\w[0][2] ),
    .Y(_10405_));
 sky130_fd_sc_hd__o21ai_4 _24553_ (.A1(net286),
    .A2(_10404_),
    .B1(_10405_),
    .Y(_00022_));
 sky130_fd_sc_hd__mux4_2 _24554_ (.A0(\w[18][3] ),
    .A1(\w[16][3] ),
    .A2(\w[22][3] ),
    .A3(\w[20][3] ),
    .S0(net365),
    .S1(net304),
    .X(_10406_));
 sky130_fd_sc_hd__mux4_2 _24555_ (.A0(\w[26][3] ),
    .A1(\w[24][3] ),
    .A2(\w[30][3] ),
    .A3(\w[28][3] ),
    .S0(net365),
    .S1(net304),
    .X(_10407_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_470 ();
 sky130_fd_sc_hd__mux4_2 _24557_ (.A0(\w[2][3] ),
    .A1(\w[0][3] ),
    .A2(\w[6][3] ),
    .A3(\w[4][3] ),
    .S0(net365),
    .S1(net304),
    .X(_10409_));
 sky130_fd_sc_hd__mux4_2 _24558_ (.A0(\w[10][3] ),
    .A1(\w[8][3] ),
    .A2(\w[14][3] ),
    .A3(\w[12][3] ),
    .S0(net365),
    .S1(net304),
    .X(_10410_));
 sky130_fd_sc_hd__mux4_2 _24559_ (.A0(_10406_),
    .A1(_10407_),
    .A2(_10409_),
    .A3(_10410_),
    .S0(net325),
    .S1(_10352_),
    .X(_10411_));
 sky130_fd_sc_hd__mux4_2 _24560_ (.A0(\w[50][3] ),
    .A1(\w[48][3] ),
    .A2(\w[54][3] ),
    .A3(\w[52][3] ),
    .S0(net366),
    .S1(net304),
    .X(_10412_));
 sky130_fd_sc_hd__mux4_2 _24561_ (.A0(\w[58][3] ),
    .A1(\w[56][3] ),
    .A2(\w[62][3] ),
    .A3(\w[60][3] ),
    .S0(net366),
    .S1(net304),
    .X(_10413_));
 sky130_fd_sc_hd__mux4_2 _24562_ (.A0(\w[34][3] ),
    .A1(\w[32][3] ),
    .A2(\w[38][3] ),
    .A3(\w[36][3] ),
    .S0(net366),
    .S1(net304),
    .X(_10414_));
 sky130_fd_sc_hd__mux4_2 _24563_ (.A0(\w[42][3] ),
    .A1(\w[40][3] ),
    .A2(\w[46][3] ),
    .A3(\w[44][3] ),
    .S0(net366),
    .S1(net304),
    .X(_10415_));
 sky130_fd_sc_hd__mux4_2 _24564_ (.A0(_10412_),
    .A1(_10413_),
    .A2(_10414_),
    .A3(_10415_),
    .S0(net325),
    .S1(_10352_),
    .X(_10416_));
 sky130_fd_sc_hd__mux2i_2 _24565_ (.A0(_10411_),
    .A1(_10416_),
    .S(net291),
    .Y(_10417_));
 sky130_fd_sc_hd__nand2_2 _24566_ (.A(reset_hash),
    .B(\w[0][3] ),
    .Y(_10418_));
 sky130_fd_sc_hd__o21ai_4 _24567_ (.A1(net286),
    .A2(_10417_),
    .B1(_10418_),
    .Y(_00025_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_469 ();
 sky130_fd_sc_hd__mux4_2 _24569_ (.A0(\w[18][4] ),
    .A1(\w[16][4] ),
    .A2(\w[22][4] ),
    .A3(\w[20][4] ),
    .S0(net368),
    .S1(net305),
    .X(_10420_));
 sky130_fd_sc_hd__mux4_2 _24570_ (.A0(\w[26][4] ),
    .A1(\w[24][4] ),
    .A2(\w[30][4] ),
    .A3(\w[28][4] ),
    .S0(net368),
    .S1(net305),
    .X(_10421_));
 sky130_fd_sc_hd__mux4_2 _24571_ (.A0(\w[2][4] ),
    .A1(\w[0][4] ),
    .A2(\w[6][4] ),
    .A3(\w[4][4] ),
    .S0(net368),
    .S1(net305),
    .X(_10422_));
 sky130_fd_sc_hd__mux4_2 _24572_ (.A0(\w[10][4] ),
    .A1(\w[8][4] ),
    .A2(\w[14][4] ),
    .A3(\w[12][4] ),
    .S0(net368),
    .S1(net305),
    .X(_10423_));
 sky130_fd_sc_hd__mux4_2 _24573_ (.A0(_10420_),
    .A1(_10421_),
    .A2(_10422_),
    .A3(_10423_),
    .S0(net322),
    .S1(net313),
    .X(_10424_));
 sky130_fd_sc_hd__mux4_2 _24574_ (.A0(\w[50][4] ),
    .A1(\w[48][4] ),
    .A2(\w[54][4] ),
    .A3(\w[52][4] ),
    .S0(net365),
    .S1(net305),
    .X(_10425_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_468 ();
 sky130_fd_sc_hd__mux4_2 _24576_ (.A0(\w[58][4] ),
    .A1(\w[56][4] ),
    .A2(\w[62][4] ),
    .A3(\w[60][4] ),
    .S0(net365),
    .S1(net305),
    .X(_10427_));
 sky130_fd_sc_hd__mux4_2 _24577_ (.A0(\w[34][4] ),
    .A1(\w[32][4] ),
    .A2(\w[38][4] ),
    .A3(\w[36][4] ),
    .S0(net365),
    .S1(net305),
    .X(_10428_));
 sky130_fd_sc_hd__mux4_2 _24578_ (.A0(\w[42][4] ),
    .A1(\w[40][4] ),
    .A2(\w[46][4] ),
    .A3(\w[44][4] ),
    .S0(net365),
    .S1(net305),
    .X(_10429_));
 sky130_fd_sc_hd__mux4_2 _24579_ (.A0(_10425_),
    .A1(_10427_),
    .A2(_10428_),
    .A3(_10429_),
    .S0(net323),
    .S1(net314),
    .X(_10430_));
 sky130_fd_sc_hd__mux2i_1 _24580_ (.A0(_10424_),
    .A1(_10430_),
    .S(net288),
    .Y(_10431_));
 sky130_fd_sc_hd__nand2_2 _24581_ (.A(reset_hash),
    .B(\w[0][4] ),
    .Y(_10432_));
 sky130_fd_sc_hd__o21ai_4 _24582_ (.A1(net286),
    .A2(_10431_),
    .B1(_10432_),
    .Y(_00026_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_467 ();
 sky130_fd_sc_hd__mux4_2 _24584_ (.A0(\w[18][5] ),
    .A1(\w[16][5] ),
    .A2(\w[22][5] ),
    .A3(\w[20][5] ),
    .S0(net365),
    .S1(net305),
    .X(_10434_));
 sky130_fd_sc_hd__mux4_2 _24585_ (.A0(\w[26][5] ),
    .A1(\w[24][5] ),
    .A2(\w[30][5] ),
    .A3(\w[28][5] ),
    .S0(net365),
    .S1(net305),
    .X(_10435_));
 sky130_fd_sc_hd__mux4_2 _24586_ (.A0(\w[2][5] ),
    .A1(\w[0][5] ),
    .A2(\w[6][5] ),
    .A3(\w[4][5] ),
    .S0(net365),
    .S1(net305),
    .X(_10436_));
 sky130_fd_sc_hd__mux4_2 _24587_ (.A0(\w[10][5] ),
    .A1(\w[8][5] ),
    .A2(\w[14][5] ),
    .A3(\w[12][5] ),
    .S0(net365),
    .S1(net305),
    .X(_10437_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_466 ();
 sky130_fd_sc_hd__mux4_2 _24589_ (.A0(_10434_),
    .A1(_10435_),
    .A2(_10436_),
    .A3(_10437_),
    .S0(net323),
    .S1(net314),
    .X(_10439_));
 sky130_fd_sc_hd__mux4_2 _24590_ (.A0(\w[50][5] ),
    .A1(\w[48][5] ),
    .A2(\w[54][5] ),
    .A3(\w[52][5] ),
    .S0(net365),
    .S1(net306),
    .X(_10440_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_465 ();
 sky130_fd_sc_hd__mux4_2 _24592_ (.A0(\w[58][5] ),
    .A1(\w[56][5] ),
    .A2(\w[62][5] ),
    .A3(\w[60][5] ),
    .S0(net365),
    .S1(net306),
    .X(_10442_));
 sky130_fd_sc_hd__mux4_2 _24593_ (.A0(\w[34][5] ),
    .A1(\w[32][5] ),
    .A2(\w[38][5] ),
    .A3(\w[36][5] ),
    .S0(net365),
    .S1(net306),
    .X(_10443_));
 sky130_fd_sc_hd__mux4_2 _24594_ (.A0(\w[42][5] ),
    .A1(\w[40][5] ),
    .A2(\w[46][5] ),
    .A3(\w[44][5] ),
    .S0(net365),
    .S1(net306),
    .X(_10444_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_464 ();
 sky130_fd_sc_hd__mux4_2 _24596_ (.A0(_10440_),
    .A1(_10442_),
    .A2(_10443_),
    .A3(_10444_),
    .S0(net323),
    .S1(net314),
    .X(_10446_));
 sky130_fd_sc_hd__mux2i_1 _24597_ (.A0(_10439_),
    .A1(_10446_),
    .S(net288),
    .Y(_10447_));
 sky130_fd_sc_hd__nand2_2 _24598_ (.A(reset_hash),
    .B(\w[0][5] ),
    .Y(_10448_));
 sky130_fd_sc_hd__o21ai_4 _24599_ (.A1(net286),
    .A2(_10447_),
    .B1(_10448_),
    .Y(_00027_));
 sky130_fd_sc_hd__mux4_2 _24600_ (.A0(\w[18][6] ),
    .A1(\w[16][6] ),
    .A2(\w[22][6] ),
    .A3(\w[20][6] ),
    .S0(net365),
    .S1(net304),
    .X(_10449_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_463 ();
 sky130_fd_sc_hd__mux4_2 _24602_ (.A0(\w[26][6] ),
    .A1(\w[24][6] ),
    .A2(\w[30][6] ),
    .A3(\w[28][6] ),
    .S0(net365),
    .S1(net304),
    .X(_10451_));
 sky130_fd_sc_hd__mux4_2 _24603_ (.A0(\w[2][6] ),
    .A1(\w[0][6] ),
    .A2(\w[6][6] ),
    .A3(\w[4][6] ),
    .S0(net365),
    .S1(net304),
    .X(_10452_));
 sky130_fd_sc_hd__mux4_2 _24604_ (.A0(\w[10][6] ),
    .A1(\w[8][6] ),
    .A2(\w[14][6] ),
    .A3(\w[12][6] ),
    .S0(net365),
    .S1(net304),
    .X(_10453_));
 sky130_fd_sc_hd__mux4_2 _24605_ (.A0(_10449_),
    .A1(_10451_),
    .A2(_10452_),
    .A3(_10453_),
    .S0(net323),
    .S1(net314),
    .X(_10454_));
 sky130_fd_sc_hd__mux4_2 _24606_ (.A0(\w[50][6] ),
    .A1(\w[48][6] ),
    .A2(\w[54][6] ),
    .A3(\w[52][6] ),
    .S0(net366),
    .S1(net304),
    .X(_10455_));
 sky130_fd_sc_hd__mux4_2 _24607_ (.A0(\w[58][6] ),
    .A1(\w[56][6] ),
    .A2(\w[62][6] ),
    .A3(\w[60][6] ),
    .S0(net366),
    .S1(net304),
    .X(_10456_));
 sky130_fd_sc_hd__mux4_2 _24608_ (.A0(\w[34][6] ),
    .A1(\w[32][6] ),
    .A2(\w[38][6] ),
    .A3(\w[36][6] ),
    .S0(net366),
    .S1(net304),
    .X(_10457_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_462 ();
 sky130_fd_sc_hd__mux4_2 _24610_ (.A0(\w[42][6] ),
    .A1(\w[40][6] ),
    .A2(\w[46][6] ),
    .A3(\w[44][6] ),
    .S0(net366),
    .S1(net304),
    .X(_10459_));
 sky130_fd_sc_hd__mux4_2 _24611_ (.A0(_10455_),
    .A1(_10456_),
    .A2(_10457_),
    .A3(_10459_),
    .S0(net323),
    .S1(net314),
    .X(_10460_));
 sky130_fd_sc_hd__mux2i_1 _24612_ (.A0(_10454_),
    .A1(_10460_),
    .S(net288),
    .Y(_10461_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_461 ();
 sky130_fd_sc_hd__nand2_2 _24614_ (.A(reset_hash),
    .B(\w[0][6] ),
    .Y(_10463_));
 sky130_fd_sc_hd__o21ai_4 _24615_ (.A1(net286),
    .A2(_10461_),
    .B1(_10463_),
    .Y(_00028_));
 sky130_fd_sc_hd__mux4_2 _24616_ (.A0(\w[18][7] ),
    .A1(\w[16][7] ),
    .A2(\w[22][7] ),
    .A3(\w[20][7] ),
    .S0(net368),
    .S1(net305),
    .X(_10464_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_460 ();
 sky130_fd_sc_hd__mux4_2 _24618_ (.A0(\w[26][7] ),
    .A1(\w[24][7] ),
    .A2(\w[30][7] ),
    .A3(\w[28][7] ),
    .S0(net368),
    .S1(net305),
    .X(_10466_));
 sky130_fd_sc_hd__mux4_2 _24619_ (.A0(\w[2][7] ),
    .A1(\w[0][7] ),
    .A2(\w[6][7] ),
    .A3(\w[4][7] ),
    .S0(net368),
    .S1(net305),
    .X(_10467_));
 sky130_fd_sc_hd__mux4_2 _24620_ (.A0(\w[10][7] ),
    .A1(\w[8][7] ),
    .A2(\w[14][7] ),
    .A3(\w[12][7] ),
    .S0(net368),
    .S1(net305),
    .X(_10468_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_459 ();
 sky130_fd_sc_hd__mux4_2 _24622_ (.A0(_10464_),
    .A1(_10466_),
    .A2(_10467_),
    .A3(_10468_),
    .S0(net322),
    .S1(net313),
    .X(_10470_));
 sky130_fd_sc_hd__mux4_2 _24623_ (.A0(\w[50][7] ),
    .A1(\w[48][7] ),
    .A2(\w[54][7] ),
    .A3(\w[52][7] ),
    .S0(net365),
    .S1(net304),
    .X(_10471_));
 sky130_fd_sc_hd__mux4_2 _24624_ (.A0(\w[58][7] ),
    .A1(\w[56][7] ),
    .A2(\w[62][7] ),
    .A3(\w[60][7] ),
    .S0(net365),
    .S1(net304),
    .X(_10472_));
 sky130_fd_sc_hd__mux4_2 _24625_ (.A0(\w[34][7] ),
    .A1(\w[32][7] ),
    .A2(\w[38][7] ),
    .A3(\w[36][7] ),
    .S0(net365),
    .S1(net304),
    .X(_10473_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_458 ();
 sky130_fd_sc_hd__mux4_2 _24627_ (.A0(\w[42][7] ),
    .A1(\w[40][7] ),
    .A2(\w[46][7] ),
    .A3(\w[44][7] ),
    .S0(net365),
    .S1(net304),
    .X(_10475_));
 sky130_fd_sc_hd__mux4_2 _24628_ (.A0(_10471_),
    .A1(_10472_),
    .A2(_10473_),
    .A3(_10475_),
    .S0(net323),
    .S1(net314),
    .X(_10476_));
 sky130_fd_sc_hd__mux2i_1 _24629_ (.A0(_10470_),
    .A1(_10476_),
    .S(net288),
    .Y(_10477_));
 sky130_fd_sc_hd__nand2_2 _24630_ (.A(net348),
    .B(\w[0][7] ),
    .Y(_10478_));
 sky130_fd_sc_hd__o21ai_4 _24631_ (.A1(net286),
    .A2(_10477_),
    .B1(_10478_),
    .Y(_00029_));
 sky130_fd_sc_hd__mux4_2 _24632_ (.A0(\w[18][8] ),
    .A1(\w[16][8] ),
    .A2(\w[22][8] ),
    .A3(\w[20][8] ),
    .S0(net371),
    .S1(net307),
    .X(_10479_));
 sky130_fd_sc_hd__mux4_2 _24633_ (.A0(\w[26][8] ),
    .A1(\w[24][8] ),
    .A2(\w[30][8] ),
    .A3(\w[28][8] ),
    .S0(net371),
    .S1(net307),
    .X(_10480_));
 sky130_fd_sc_hd__mux4_2 _24634_ (.A0(\w[2][8] ),
    .A1(\w[0][8] ),
    .A2(\w[6][8] ),
    .A3(\w[4][8] ),
    .S0(net371),
    .S1(net307),
    .X(_10481_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_457 ();
 sky130_fd_sc_hd__mux4_2 _24636_ (.A0(\w[10][8] ),
    .A1(\w[8][8] ),
    .A2(\w[14][8] ),
    .A3(\w[12][8] ),
    .S0(net371),
    .S1(net307),
    .X(_10483_));
 sky130_fd_sc_hd__mux4_2 _24637_ (.A0(_10479_),
    .A1(_10480_),
    .A2(_10481_),
    .A3(_10483_),
    .S0(net321),
    .S1(net317),
    .X(_10484_));
 sky130_fd_sc_hd__mux4_2 _24638_ (.A0(\w[50][8] ),
    .A1(\w[48][8] ),
    .A2(\w[54][8] ),
    .A3(\w[52][8] ),
    .S0(net368),
    .S1(net305),
    .X(_10485_));
 sky130_fd_sc_hd__mux4_2 _24639_ (.A0(\w[58][8] ),
    .A1(\w[56][8] ),
    .A2(\w[62][8] ),
    .A3(\w[60][8] ),
    .S0(net368),
    .S1(net305),
    .X(_10486_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_456 ();
 sky130_fd_sc_hd__mux4_2 _24641_ (.A0(\w[34][8] ),
    .A1(\w[32][8] ),
    .A2(\w[38][8] ),
    .A3(\w[36][8] ),
    .S0(net368),
    .S1(net305),
    .X(_10488_));
 sky130_fd_sc_hd__mux4_2 _24642_ (.A0(\w[42][8] ),
    .A1(\w[40][8] ),
    .A2(\w[46][8] ),
    .A3(\w[44][8] ),
    .S0(net368),
    .S1(net305),
    .X(_10489_));
 sky130_fd_sc_hd__mux4_2 _24643_ (.A0(_10485_),
    .A1(_10486_),
    .A2(_10488_),
    .A3(_10489_),
    .S0(net324),
    .S1(net315),
    .X(_10490_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_454 ();
 sky130_fd_sc_hd__mux2i_1 _24646_ (.A0(_10484_),
    .A1(_10490_),
    .S(net289),
    .Y(_10493_));
 sky130_fd_sc_hd__nand2_1 _24647_ (.A(net348),
    .B(\w[0][8] ),
    .Y(_10494_));
 sky130_fd_sc_hd__o21ai_1 _24648_ (.A1(net286),
    .A2(_10493_),
    .B1(_10494_),
    .Y(_00030_));
 sky130_fd_sc_hd__mux4_2 _24649_ (.A0(\w[18][9] ),
    .A1(\w[16][9] ),
    .A2(\w[22][9] ),
    .A3(\w[20][9] ),
    .S0(net371),
    .S1(net307),
    .X(_10495_));
 sky130_fd_sc_hd__mux4_2 _24650_ (.A0(\w[26][9] ),
    .A1(\w[24][9] ),
    .A2(\w[30][9] ),
    .A3(\w[28][9] ),
    .S0(net371),
    .S1(net307),
    .X(_10496_));
 sky130_fd_sc_hd__mux4_2 _24651_ (.A0(\w[2][9] ),
    .A1(\w[0][9] ),
    .A2(\w[6][9] ),
    .A3(\w[4][9] ),
    .S0(net371),
    .S1(net307),
    .X(_10497_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_453 ();
 sky130_fd_sc_hd__mux4_2 _24653_ (.A0(\w[10][9] ),
    .A1(\w[8][9] ),
    .A2(\w[14][9] ),
    .A3(\w[12][9] ),
    .S0(net371),
    .S1(net307),
    .X(_10499_));
 sky130_fd_sc_hd__mux4_2 _24654_ (.A0(_10495_),
    .A1(_10496_),
    .A2(_10497_),
    .A3(_10499_),
    .S0(net320),
    .S1(net316),
    .X(_10500_));
 sky130_fd_sc_hd__mux4_2 _24655_ (.A0(\w[50][9] ),
    .A1(\w[48][9] ),
    .A2(\w[54][9] ),
    .A3(\w[52][9] ),
    .S0(net370),
    .S1(net306),
    .X(_10501_));
 sky130_fd_sc_hd__mux4_2 _24656_ (.A0(\w[58][9] ),
    .A1(\w[56][9] ),
    .A2(\w[62][9] ),
    .A3(\w[60][9] ),
    .S0(net370),
    .S1(net306),
    .X(_10502_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_452 ();
 sky130_fd_sc_hd__mux4_2 _24658_ (.A0(\w[34][9] ),
    .A1(\w[32][9] ),
    .A2(\w[38][9] ),
    .A3(\w[36][9] ),
    .S0(net370),
    .S1(net306),
    .X(_10504_));
 sky130_fd_sc_hd__mux4_2 _24659_ (.A0(\w[42][9] ),
    .A1(\w[40][9] ),
    .A2(\w[46][9] ),
    .A3(\w[44][9] ),
    .S0(net370),
    .S1(net306),
    .X(_10505_));
 sky130_fd_sc_hd__mux4_2 _24660_ (.A0(_10501_),
    .A1(_10502_),
    .A2(_10504_),
    .A3(_10505_),
    .S0(net324),
    .S1(net315),
    .X(_10506_));
 sky130_fd_sc_hd__mux2i_1 _24661_ (.A0(_10500_),
    .A1(_10506_),
    .S(net290),
    .Y(_10507_));
 sky130_fd_sc_hd__nand2_1 _24662_ (.A(net348),
    .B(\w[0][9] ),
    .Y(_10508_));
 sky130_fd_sc_hd__o21ai_0 _24663_ (.A1(net287),
    .A2(_10507_),
    .B1(_10508_),
    .Y(_00031_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_451 ();
 sky130_fd_sc_hd__mux4_2 _24665_ (.A0(\w[18][10] ),
    .A1(\w[16][10] ),
    .A2(\w[22][10] ),
    .A3(\w[20][10] ),
    .S0(net371),
    .S1(net307),
    .X(_10510_));
 sky130_fd_sc_hd__mux4_2 _24666_ (.A0(\w[26][10] ),
    .A1(\w[24][10] ),
    .A2(\w[30][10] ),
    .A3(\w[28][10] ),
    .S0(net371),
    .S1(net307),
    .X(_10511_));
 sky130_fd_sc_hd__mux4_2 _24667_ (.A0(\w[2][10] ),
    .A1(\w[0][10] ),
    .A2(\w[6][10] ),
    .A3(\w[4][10] ),
    .S0(net371),
    .S1(net307),
    .X(_10512_));
 sky130_fd_sc_hd__mux4_2 _24668_ (.A0(\w[10][10] ),
    .A1(\w[8][10] ),
    .A2(\w[14][10] ),
    .A3(\w[12][10] ),
    .S0(net371),
    .S1(net307),
    .X(_10513_));
 sky130_fd_sc_hd__mux4_2 _24669_ (.A0(_10510_),
    .A1(_10511_),
    .A2(_10512_),
    .A3(_10513_),
    .S0(net320),
    .S1(net318),
    .X(_10514_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_450 ();
 sky130_fd_sc_hd__mux4_2 _24671_ (.A0(\w[50][10] ),
    .A1(\w[48][10] ),
    .A2(\w[54][10] ),
    .A3(\w[52][10] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10516_));
 sky130_fd_sc_hd__mux4_2 _24672_ (.A0(\w[58][10] ),
    .A1(\w[56][10] ),
    .A2(\w[62][10] ),
    .A3(\w[60][10] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10517_));
 sky130_fd_sc_hd__mux4_2 _24673_ (.A0(\w[34][10] ),
    .A1(\w[32][10] ),
    .A2(\w[38][10] ),
    .A3(\w[36][10] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10518_));
 sky130_fd_sc_hd__mux4_2 _24674_ (.A0(\w[42][10] ),
    .A1(\w[40][10] ),
    .A2(\w[46][10] ),
    .A3(\w[44][10] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10519_));
 sky130_fd_sc_hd__mux4_2 _24675_ (.A0(_10516_),
    .A1(_10517_),
    .A2(_10518_),
    .A3(_10519_),
    .S0(_10348_),
    .S1(net317),
    .X(_10520_));
 sky130_fd_sc_hd__mux2i_1 _24676_ (.A0(_10514_),
    .A1(_10520_),
    .S(_10373_),
    .Y(_10521_));
 sky130_fd_sc_hd__nand2_1 _24677_ (.A(net348),
    .B(\w[0][10] ),
    .Y(_10522_));
 sky130_fd_sc_hd__o21ai_0 _24678_ (.A1(net287),
    .A2(_10521_),
    .B1(_10522_),
    .Y(_00001_));
 sky130_fd_sc_hd__mux4_2 _24679_ (.A0(\w[18][11] ),
    .A1(\w[16][11] ),
    .A2(\w[22][11] ),
    .A3(\w[20][11] ),
    .S0(net369),
    .S1(net307),
    .X(_10523_));
 sky130_fd_sc_hd__mux4_2 _24680_ (.A0(\w[26][11] ),
    .A1(\w[24][11] ),
    .A2(\w[30][11] ),
    .A3(\w[28][11] ),
    .S0(net369),
    .S1(net307),
    .X(_10524_));
 sky130_fd_sc_hd__mux4_2 _24681_ (.A0(\w[2][11] ),
    .A1(\w[0][11] ),
    .A2(\w[6][11] ),
    .A3(\w[4][11] ),
    .S0(net369),
    .S1(net307),
    .X(_10525_));
 sky130_fd_sc_hd__mux4_2 _24682_ (.A0(\w[10][11] ),
    .A1(\w[8][11] ),
    .A2(\w[14][11] ),
    .A3(\w[12][11] ),
    .S0(net369),
    .S1(net307),
    .X(_10526_));
 sky130_fd_sc_hd__mux4_2 _24683_ (.A0(_10523_),
    .A1(_10524_),
    .A2(_10525_),
    .A3(_10526_),
    .S0(net321),
    .S1(net317),
    .X(_10527_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_449 ();
 sky130_fd_sc_hd__mux4_2 _24685_ (.A0(\w[50][11] ),
    .A1(\w[48][11] ),
    .A2(\w[54][11] ),
    .A3(\w[52][11] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10529_));
 sky130_fd_sc_hd__mux4_2 _24686_ (.A0(\w[58][11] ),
    .A1(\w[56][11] ),
    .A2(\w[62][11] ),
    .A3(\w[60][11] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10530_));
 sky130_fd_sc_hd__mux4_2 _24687_ (.A0(\w[34][11] ),
    .A1(\w[32][11] ),
    .A2(\w[38][11] ),
    .A3(\w[36][11] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10531_));
 sky130_fd_sc_hd__mux4_2 _24688_ (.A0(\w[42][11] ),
    .A1(\w[40][11] ),
    .A2(\w[46][11] ),
    .A3(\w[44][11] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10532_));
 sky130_fd_sc_hd__mux4_2 _24689_ (.A0(_10529_),
    .A1(_10530_),
    .A2(_10531_),
    .A3(_10532_),
    .S0(net325),
    .S1(_10352_),
    .X(_10533_));
 sky130_fd_sc_hd__mux2i_1 _24690_ (.A0(_10527_),
    .A1(_10533_),
    .S(net289),
    .Y(_10534_));
 sky130_fd_sc_hd__nand2_2 _24691_ (.A(net348),
    .B(\w[0][11] ),
    .Y(_10535_));
 sky130_fd_sc_hd__o21ai_4 _24692_ (.A1(net286),
    .A2(_10534_),
    .B1(_10535_),
    .Y(_00002_));
 sky130_fd_sc_hd__mux4_2 _24693_ (.A0(\w[18][12] ),
    .A1(\w[16][12] ),
    .A2(\w[22][12] ),
    .A3(\w[20][12] ),
    .S0(net368),
    .S1(net305),
    .X(_10536_));
 sky130_fd_sc_hd__mux4_2 _24694_ (.A0(\w[26][12] ),
    .A1(\w[24][12] ),
    .A2(\w[30][12] ),
    .A3(\w[28][12] ),
    .S0(net368),
    .S1(net305),
    .X(_10537_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_448 ();
 sky130_fd_sc_hd__mux4_2 _24696_ (.A0(\w[2][12] ),
    .A1(\w[0][12] ),
    .A2(\w[6][12] ),
    .A3(\w[4][12] ),
    .S0(net368),
    .S1(net305),
    .X(_10539_));
 sky130_fd_sc_hd__mux4_2 _24697_ (.A0(\w[10][12] ),
    .A1(\w[8][12] ),
    .A2(\w[14][12] ),
    .A3(\w[12][12] ),
    .S0(net368),
    .S1(net305),
    .X(_10540_));
 sky130_fd_sc_hd__mux4_2 _24698_ (.A0(_10536_),
    .A1(_10537_),
    .A2(_10539_),
    .A3(_10540_),
    .S0(net322),
    .S1(net313),
    .X(_10541_));
 sky130_fd_sc_hd__mux4_2 _24699_ (.A0(\w[50][12] ),
    .A1(\w[48][12] ),
    .A2(\w[54][12] ),
    .A3(\w[52][12] ),
    .S0(net366),
    .S1(net304),
    .X(_10542_));
 sky130_fd_sc_hd__mux4_2 _24700_ (.A0(\w[58][12] ),
    .A1(\w[56][12] ),
    .A2(\w[62][12] ),
    .A3(\w[60][12] ),
    .S0(net366),
    .S1(net304),
    .X(_10543_));
 sky130_fd_sc_hd__mux4_2 _24701_ (.A0(\w[34][12] ),
    .A1(\w[32][12] ),
    .A2(\w[38][12] ),
    .A3(\w[36][12] ),
    .S0(net366),
    .S1(net304),
    .X(_10544_));
 sky130_fd_sc_hd__mux4_2 _24702_ (.A0(\w[42][12] ),
    .A1(\w[40][12] ),
    .A2(\w[46][12] ),
    .A3(\w[44][12] ),
    .S0(net366),
    .S1(net306),
    .X(_10545_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_447 ();
 sky130_fd_sc_hd__mux4_2 _24704_ (.A0(_10542_),
    .A1(_10543_),
    .A2(_10544_),
    .A3(_10545_),
    .S0(net323),
    .S1(net314),
    .X(_10547_));
 sky130_fd_sc_hd__mux2i_1 _24705_ (.A0(_10541_),
    .A1(_10547_),
    .S(net288),
    .Y(_10548_));
 sky130_fd_sc_hd__nand2_2 _24706_ (.A(net348),
    .B(\w[0][12] ),
    .Y(_10549_));
 sky130_fd_sc_hd__o21ai_4 _24707_ (.A1(net286),
    .A2(_10548_),
    .B1(_10549_),
    .Y(_00003_));
 sky130_fd_sc_hd__mux4_2 _24708_ (.A0(\w[18][13] ),
    .A1(\w[16][13] ),
    .A2(\w[22][13] ),
    .A3(\w[20][13] ),
    .S0(net367),
    .S1(net305),
    .X(_10550_));
 sky130_fd_sc_hd__mux4_2 _24709_ (.A0(\w[26][13] ),
    .A1(\w[24][13] ),
    .A2(\w[30][13] ),
    .A3(\w[28][13] ),
    .S0(net367),
    .S1(net305),
    .X(_10551_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_446 ();
 sky130_fd_sc_hd__mux4_2 _24711_ (.A0(\w[2][13] ),
    .A1(\w[0][13] ),
    .A2(\w[6][13] ),
    .A3(\w[4][13] ),
    .S0(net367),
    .S1(net305),
    .X(_10553_));
 sky130_fd_sc_hd__mux4_2 _24712_ (.A0(\w[10][13] ),
    .A1(\w[8][13] ),
    .A2(\w[14][13] ),
    .A3(\w[12][13] ),
    .S0(net367),
    .S1(net305),
    .X(_10554_));
 sky130_fd_sc_hd__mux4_2 _24713_ (.A0(_10550_),
    .A1(_10551_),
    .A2(_10553_),
    .A3(_10554_),
    .S0(net324),
    .S1(net315),
    .X(_10555_));
 sky130_fd_sc_hd__mux4_2 _24714_ (.A0(\w[50][13] ),
    .A1(\w[48][13] ),
    .A2(\w[54][13] ),
    .A3(\w[52][13] ),
    .S0(net366),
    .S1(net304),
    .X(_10556_));
 sky130_fd_sc_hd__mux4_2 _24715_ (.A0(\w[58][13] ),
    .A1(\w[56][13] ),
    .A2(\w[62][13] ),
    .A3(\w[60][13] ),
    .S0(net366),
    .S1(net304),
    .X(_10557_));
 sky130_fd_sc_hd__mux4_2 _24716_ (.A0(\w[34][13] ),
    .A1(\w[32][13] ),
    .A2(\w[38][13] ),
    .A3(\w[36][13] ),
    .S0(net366),
    .S1(net304),
    .X(_10558_));
 sky130_fd_sc_hd__mux4_2 _24717_ (.A0(\w[42][13] ),
    .A1(\w[40][13] ),
    .A2(\w[46][13] ),
    .A3(\w[44][13] ),
    .S0(net366),
    .S1(net304),
    .X(_10559_));
 sky130_fd_sc_hd__mux4_2 _24718_ (.A0(_10556_),
    .A1(_10557_),
    .A2(_10558_),
    .A3(_10559_),
    .S0(net323),
    .S1(net314),
    .X(_10560_));
 sky130_fd_sc_hd__mux2i_1 _24719_ (.A0(_10555_),
    .A1(_10560_),
    .S(net288),
    .Y(_10561_));
 sky130_fd_sc_hd__nand2_2 _24720_ (.A(net348),
    .B(\w[0][13] ),
    .Y(_10562_));
 sky130_fd_sc_hd__o21ai_4 _24721_ (.A1(net286),
    .A2(_10561_),
    .B1(_10562_),
    .Y(_00004_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_445 ();
 sky130_fd_sc_hd__mux4_2 _24723_ (.A0(\w[18][14] ),
    .A1(\w[16][14] ),
    .A2(\w[22][14] ),
    .A3(\w[20][14] ),
    .S0(net369),
    .S1(net303),
    .X(_10564_));
 sky130_fd_sc_hd__mux4_2 _24724_ (.A0(\w[26][14] ),
    .A1(\w[24][14] ),
    .A2(\w[30][14] ),
    .A3(\w[28][14] ),
    .S0(net369),
    .S1(net303),
    .X(_10565_));
 sky130_fd_sc_hd__mux4_2 _24725_ (.A0(\w[2][14] ),
    .A1(\w[0][14] ),
    .A2(\w[6][14] ),
    .A3(\w[4][14] ),
    .S0(net369),
    .S1(net303),
    .X(_10566_));
 sky130_fd_sc_hd__mux4_2 _24726_ (.A0(\w[10][14] ),
    .A1(\w[8][14] ),
    .A2(\w[14][14] ),
    .A3(\w[12][14] ),
    .S0(net369),
    .S1(net303),
    .X(_10567_));
 sky130_fd_sc_hd__mux4_2 _24727_ (.A0(_10564_),
    .A1(_10565_),
    .A2(_10566_),
    .A3(_10567_),
    .S0(net321),
    .S1(net317),
    .X(_10568_));
 sky130_fd_sc_hd__mux4_2 _24728_ (.A0(\w[50][14] ),
    .A1(\w[48][14] ),
    .A2(\w[54][14] ),
    .A3(\w[52][14] ),
    .S0(net366),
    .S1(net304),
    .X(_10569_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_444 ();
 sky130_fd_sc_hd__mux4_2 _24730_ (.A0(\w[58][14] ),
    .A1(\w[56][14] ),
    .A2(\w[62][14] ),
    .A3(\w[60][14] ),
    .S0(net366),
    .S1(net306),
    .X(_10571_));
 sky130_fd_sc_hd__mux4_2 _24731_ (.A0(\w[34][14] ),
    .A1(\w[32][14] ),
    .A2(\w[38][14] ),
    .A3(\w[36][14] ),
    .S0(net370),
    .S1(net306),
    .X(_10572_));
 sky130_fd_sc_hd__mux4_2 _24732_ (.A0(\w[42][14] ),
    .A1(\w[40][14] ),
    .A2(\w[46][14] ),
    .A3(\w[44][14] ),
    .S0(net366),
    .S1(net306),
    .X(_10573_));
 sky130_fd_sc_hd__mux4_2 _24733_ (.A0(_10569_),
    .A1(_10571_),
    .A2(_10572_),
    .A3(_10573_),
    .S0(net324),
    .S1(net314),
    .X(_10574_));
 sky130_fd_sc_hd__mux2i_1 _24734_ (.A0(_10568_),
    .A1(_10574_),
    .S(net288),
    .Y(_10575_));
 sky130_fd_sc_hd__nand2_1 _24735_ (.A(net348),
    .B(\w[0][14] ),
    .Y(_10576_));
 sky130_fd_sc_hd__o21ai_2 _24736_ (.A1(net286),
    .A2(_10575_),
    .B1(_10576_),
    .Y(_00005_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_443 ();
 sky130_fd_sc_hd__mux4_2 _24738_ (.A0(\w[18][15] ),
    .A1(\w[16][15] ),
    .A2(\w[22][15] ),
    .A3(\w[20][15] ),
    .S0(net365),
    .S1(net306),
    .X(_10578_));
 sky130_fd_sc_hd__mux4_2 _24739_ (.A0(\w[26][15] ),
    .A1(\w[24][15] ),
    .A2(\w[30][15] ),
    .A3(\w[28][15] ),
    .S0(net365),
    .S1(net306),
    .X(_10579_));
 sky130_fd_sc_hd__mux4_2 _24740_ (.A0(\w[2][15] ),
    .A1(\w[0][15] ),
    .A2(\w[6][15] ),
    .A3(\w[4][15] ),
    .S0(net365),
    .S1(net306),
    .X(_10580_));
 sky130_fd_sc_hd__mux4_2 _24741_ (.A0(\w[10][15] ),
    .A1(\w[8][15] ),
    .A2(\w[14][15] ),
    .A3(\w[12][15] ),
    .S0(net365),
    .S1(net306),
    .X(_10581_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_442 ();
 sky130_fd_sc_hd__mux4_2 _24743_ (.A0(_10578_),
    .A1(_10579_),
    .A2(_10580_),
    .A3(_10581_),
    .S0(net323),
    .S1(net314),
    .X(_10583_));
 sky130_fd_sc_hd__mux4_2 _24744_ (.A0(\w[50][15] ),
    .A1(\w[48][15] ),
    .A2(\w[54][15] ),
    .A3(\w[52][15] ),
    .S0(net365),
    .S1(net304),
    .X(_10584_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_441 ();
 sky130_fd_sc_hd__mux4_2 _24746_ (.A0(\w[58][15] ),
    .A1(\w[56][15] ),
    .A2(\w[62][15] ),
    .A3(\w[60][15] ),
    .S0(net365),
    .S1(net304),
    .X(_10586_));
 sky130_fd_sc_hd__mux4_2 _24747_ (.A0(\w[34][15] ),
    .A1(\w[32][15] ),
    .A2(\w[38][15] ),
    .A3(\w[36][15] ),
    .S0(net365),
    .S1(net304),
    .X(_10587_));
 sky130_fd_sc_hd__mux4_2 _24748_ (.A0(\w[42][15] ),
    .A1(\w[40][15] ),
    .A2(\w[46][15] ),
    .A3(\w[44][15] ),
    .S0(net365),
    .S1(net304),
    .X(_10588_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_440 ();
 sky130_fd_sc_hd__mux4_2 _24750_ (.A0(_10584_),
    .A1(_10586_),
    .A2(_10587_),
    .A3(_10588_),
    .S0(net323),
    .S1(net314),
    .X(_10590_));
 sky130_fd_sc_hd__mux2i_1 _24751_ (.A0(_10583_),
    .A1(_10590_),
    .S(net288),
    .Y(_10591_));
 sky130_fd_sc_hd__nand2_2 _24752_ (.A(reset_hash),
    .B(\w[0][15] ),
    .Y(_10592_));
 sky130_fd_sc_hd__o21ai_4 _24753_ (.A1(net286),
    .A2(_10591_),
    .B1(_10592_),
    .Y(_00006_));
 sky130_fd_sc_hd__mux4_2 _24754_ (.A0(\w[18][16] ),
    .A1(\w[16][16] ),
    .A2(\w[22][16] ),
    .A3(\w[20][16] ),
    .S0(net365),
    .S1(net304),
    .X(_10593_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_439 ();
 sky130_fd_sc_hd__mux4_2 _24756_ (.A0(\w[26][16] ),
    .A1(\w[24][16] ),
    .A2(\w[30][16] ),
    .A3(\w[28][16] ),
    .S0(net365),
    .S1(net304),
    .X(_10595_));
 sky130_fd_sc_hd__mux4_2 _24757_ (.A0(\w[2][16] ),
    .A1(\w[0][16] ),
    .A2(\w[6][16] ),
    .A3(\w[4][16] ),
    .S0(net365),
    .S1(net304),
    .X(_10596_));
 sky130_fd_sc_hd__mux4_2 _24758_ (.A0(\w[10][16] ),
    .A1(\w[8][16] ),
    .A2(\w[14][16] ),
    .A3(\w[12][16] ),
    .S0(net365),
    .S1(net304),
    .X(_10597_));
 sky130_fd_sc_hd__mux4_2 _24759_ (.A0(_10593_),
    .A1(_10595_),
    .A2(_10596_),
    .A3(_10597_),
    .S0(net323),
    .S1(net314),
    .X(_10598_));
 sky130_fd_sc_hd__mux4_2 _24760_ (.A0(\w[50][16] ),
    .A1(\w[48][16] ),
    .A2(\w[54][16] ),
    .A3(\w[52][16] ),
    .S0(net366),
    .S1(net304),
    .X(_10599_));
 sky130_fd_sc_hd__mux4_2 _24761_ (.A0(\w[58][16] ),
    .A1(\w[56][16] ),
    .A2(\w[62][16] ),
    .A3(\w[60][16] ),
    .S0(net366),
    .S1(net304),
    .X(_10600_));
 sky130_fd_sc_hd__mux4_2 _24762_ (.A0(\w[34][16] ),
    .A1(\w[32][16] ),
    .A2(\w[38][16] ),
    .A3(\w[36][16] ),
    .S0(net366),
    .S1(net304),
    .X(_10601_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_438 ();
 sky130_fd_sc_hd__mux4_2 _24764_ (.A0(\w[42][16] ),
    .A1(\w[40][16] ),
    .A2(\w[46][16] ),
    .A3(\w[44][16] ),
    .S0(net366),
    .S1(net304),
    .X(_10603_));
 sky130_fd_sc_hd__mux4_2 _24765_ (.A0(_10599_),
    .A1(_10600_),
    .A2(_10601_),
    .A3(_10603_),
    .S0(net325),
    .S1(_10352_),
    .X(_10604_));
 sky130_fd_sc_hd__mux2i_1 _24766_ (.A0(_10598_),
    .A1(_10604_),
    .S(net291),
    .Y(_10605_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_437 ();
 sky130_fd_sc_hd__nand2_4 _24768_ (.A(reset_hash),
    .B(\w[0][16] ),
    .Y(_10607_));
 sky130_fd_sc_hd__o21ai_4 _24769_ (.A1(net287),
    .A2(_10605_),
    .B1(_10607_),
    .Y(_00007_));
 sky130_fd_sc_hd__mux4_2 _24770_ (.A0(\w[18][17] ),
    .A1(\w[16][17] ),
    .A2(\w[22][17] ),
    .A3(\w[20][17] ),
    .S0(net369),
    .S1(net303),
    .X(_10608_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_436 ();
 sky130_fd_sc_hd__mux4_2 _24772_ (.A0(\w[26][17] ),
    .A1(\w[24][17] ),
    .A2(\w[30][17] ),
    .A3(\w[28][17] ),
    .S0(net369),
    .S1(net303),
    .X(_10610_));
 sky130_fd_sc_hd__mux4_2 _24773_ (.A0(\w[2][17] ),
    .A1(\w[0][17] ),
    .A2(\w[6][17] ),
    .A3(\w[4][17] ),
    .S0(net369),
    .S1(net303),
    .X(_10611_));
 sky130_fd_sc_hd__mux4_2 _24774_ (.A0(\w[10][17] ),
    .A1(\w[8][17] ),
    .A2(\w[14][17] ),
    .A3(\w[12][17] ),
    .S0(net369),
    .S1(net303),
    .X(_10612_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_435 ();
 sky130_fd_sc_hd__mux4_2 _24776_ (.A0(_10608_),
    .A1(_10610_),
    .A2(_10611_),
    .A3(_10612_),
    .S0(net321),
    .S1(net317),
    .X(_10614_));
 sky130_fd_sc_hd__mux4_2 _24777_ (.A0(\w[50][17] ),
    .A1(\w[48][17] ),
    .A2(\w[54][17] ),
    .A3(\w[52][17] ),
    .S0(net367),
    .S1(net305),
    .X(_10615_));
 sky130_fd_sc_hd__mux4_2 _24778_ (.A0(\w[58][17] ),
    .A1(\w[56][17] ),
    .A2(\w[62][17] ),
    .A3(\w[60][17] ),
    .S0(net368),
    .S1(net305),
    .X(_10616_));
 sky130_fd_sc_hd__mux4_2 _24779_ (.A0(\w[34][17] ),
    .A1(\w[32][17] ),
    .A2(\w[38][17] ),
    .A3(\w[36][17] ),
    .S0(net368),
    .S1(net305),
    .X(_10617_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_434 ();
 sky130_fd_sc_hd__mux4_2 _24781_ (.A0(\w[42][17] ),
    .A1(\w[40][17] ),
    .A2(\w[46][17] ),
    .A3(\w[44][17] ),
    .S0(net367),
    .S1(net305),
    .X(_10619_));
 sky130_fd_sc_hd__mux4_2 _24782_ (.A0(_10615_),
    .A1(_10616_),
    .A2(_10617_),
    .A3(_10619_),
    .S0(net324),
    .S1(net315),
    .X(_10620_));
 sky130_fd_sc_hd__mux2i_1 _24783_ (.A0(_10614_),
    .A1(_10620_),
    .S(net288),
    .Y(_10621_));
 sky130_fd_sc_hd__nand2_2 _24784_ (.A(net348),
    .B(\w[0][17] ),
    .Y(_10622_));
 sky130_fd_sc_hd__o21ai_4 _24785_ (.A1(net286),
    .A2(_10621_),
    .B1(_10622_),
    .Y(_00008_));
 sky130_fd_sc_hd__mux4_2 _24786_ (.A0(\w[18][18] ),
    .A1(\w[16][18] ),
    .A2(\w[22][18] ),
    .A3(\w[20][18] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_10623_));
 sky130_fd_sc_hd__mux4_2 _24787_ (.A0(\w[26][18] ),
    .A1(\w[24][18] ),
    .A2(\w[30][18] ),
    .A3(\w[28][18] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_10624_));
 sky130_fd_sc_hd__mux4_2 _24788_ (.A0(\w[2][18] ),
    .A1(\w[0][18] ),
    .A2(\w[6][18] ),
    .A3(\w[4][18] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_10625_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_433 ();
 sky130_fd_sc_hd__mux4_2 _24790_ (.A0(\w[10][18] ),
    .A1(\w[8][18] ),
    .A2(\w[14][18] ),
    .A3(\w[12][18] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_10627_));
 sky130_fd_sc_hd__mux4_2 _24791_ (.A0(_10623_),
    .A1(_10624_),
    .A2(_10625_),
    .A3(_10627_),
    .S0(_10348_),
    .S1(net318),
    .X(_10628_));
 sky130_fd_sc_hd__mux4_2 _24792_ (.A0(\w[50][18] ),
    .A1(\w[48][18] ),
    .A2(\w[54][18] ),
    .A3(\w[52][18] ),
    .S0(net370),
    .S1(_00655_),
    .X(_10629_));
 sky130_fd_sc_hd__mux4_2 _24793_ (.A0(\w[58][18] ),
    .A1(\w[56][18] ),
    .A2(\w[62][18] ),
    .A3(\w[60][18] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10630_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_432 ();
 sky130_fd_sc_hd__mux4_2 _24795_ (.A0(\w[34][18] ),
    .A1(\w[32][18] ),
    .A2(\w[38][18] ),
    .A3(\w[36][18] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10632_));
 sky130_fd_sc_hd__mux4_2 _24796_ (.A0(\w[42][18] ),
    .A1(\w[40][18] ),
    .A2(\w[46][18] ),
    .A3(\w[44][18] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10633_));
 sky130_fd_sc_hd__mux4_2 _24797_ (.A0(_10629_),
    .A1(_10630_),
    .A2(_10632_),
    .A3(_10633_),
    .S0(net325),
    .S1(net315),
    .X(_10634_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_431 ();
 sky130_fd_sc_hd__mux2i_1 _24799_ (.A0(_10628_),
    .A1(_10634_),
    .S(_10373_),
    .Y(_10636_));
 sky130_fd_sc_hd__nand2_1 _24800_ (.A(net349),
    .B(\w[0][18] ),
    .Y(_10637_));
 sky130_fd_sc_hd__o21ai_2 _24801_ (.A1(net287),
    .A2(_10636_),
    .B1(_10637_),
    .Y(_00009_));
 sky130_fd_sc_hd__mux4_2 _24802_ (.A0(\w[18][19] ),
    .A1(\w[16][19] ),
    .A2(\w[22][19] ),
    .A3(\w[20][19] ),
    .S0(net371),
    .S1(net307),
    .X(_10638_));
 sky130_fd_sc_hd__mux4_2 _24803_ (.A0(\w[26][19] ),
    .A1(\w[24][19] ),
    .A2(\w[30][19] ),
    .A3(\w[28][19] ),
    .S0(net371),
    .S1(net307),
    .X(_10639_));
 sky130_fd_sc_hd__mux4_2 _24804_ (.A0(\w[2][19] ),
    .A1(\w[0][19] ),
    .A2(\w[6][19] ),
    .A3(\w[4][19] ),
    .S0(net371),
    .S1(net307),
    .X(_10640_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_430 ();
 sky130_fd_sc_hd__mux4_2 _24806_ (.A0(\w[10][19] ),
    .A1(\w[8][19] ),
    .A2(\w[14][19] ),
    .A3(\w[12][19] ),
    .S0(net371),
    .S1(net307),
    .X(_10642_));
 sky130_fd_sc_hd__mux4_2 _24807_ (.A0(_10638_),
    .A1(_10639_),
    .A2(_10640_),
    .A3(_10642_),
    .S0(net320),
    .S1(net316),
    .X(_10643_));
 sky130_fd_sc_hd__mux4_2 _24808_ (.A0(\w[50][19] ),
    .A1(\w[48][19] ),
    .A2(\w[54][19] ),
    .A3(\w[52][19] ),
    .S0(net372),
    .S1(net306),
    .X(_10644_));
 sky130_fd_sc_hd__mux4_2 _24809_ (.A0(\w[58][19] ),
    .A1(\w[56][19] ),
    .A2(\w[62][19] ),
    .A3(\w[60][19] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10645_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_429 ();
 sky130_fd_sc_hd__mux4_2 _24811_ (.A0(\w[34][19] ),
    .A1(\w[32][19] ),
    .A2(\w[38][19] ),
    .A3(\w[36][19] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10647_));
 sky130_fd_sc_hd__mux4_2 _24812_ (.A0(\w[42][19] ),
    .A1(\w[40][19] ),
    .A2(\w[46][19] ),
    .A3(\w[44][19] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10648_));
 sky130_fd_sc_hd__mux4_2 _24813_ (.A0(_10644_),
    .A1(_10645_),
    .A2(_10647_),
    .A3(_10648_),
    .S0(_10348_),
    .S1(net317),
    .X(_10649_));
 sky130_fd_sc_hd__mux2i_1 _24814_ (.A0(_10643_),
    .A1(_10649_),
    .S(net289),
    .Y(_10650_));
 sky130_fd_sc_hd__nand2_1 _24815_ (.A(net348),
    .B(\w[0][19] ),
    .Y(_10651_));
 sky130_fd_sc_hd__o21ai_2 _24816_ (.A1(net286),
    .A2(_10650_),
    .B1(_10651_),
    .Y(_00010_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_428 ();
 sky130_fd_sc_hd__mux4_2 _24818_ (.A0(\w[18][20] ),
    .A1(\w[16][20] ),
    .A2(\w[22][20] ),
    .A3(\w[20][20] ),
    .S0(\count_hash1[1] ),
    .S1(_00655_),
    .X(_10653_));
 sky130_fd_sc_hd__mux4_2 _24819_ (.A0(\w[26][20] ),
    .A1(\w[24][20] ),
    .A2(\w[30][20] ),
    .A3(\w[28][20] ),
    .S0(net371),
    .S1(_00655_),
    .X(_10654_));
 sky130_fd_sc_hd__mux4_2 _24820_ (.A0(\w[2][20] ),
    .A1(\w[0][20] ),
    .A2(\w[6][20] ),
    .A3(\w[4][20] ),
    .S0(net371),
    .S1(_00655_),
    .X(_10655_));
 sky130_fd_sc_hd__mux4_2 _24821_ (.A0(\w[10][20] ),
    .A1(\w[8][20] ),
    .A2(\w[14][20] ),
    .A3(\w[12][20] ),
    .S0(net371),
    .S1(_00655_),
    .X(_10656_));
 sky130_fd_sc_hd__mux4_2 _24822_ (.A0(_10653_),
    .A1(_10654_),
    .A2(_10655_),
    .A3(_10656_),
    .S0(net320),
    .S1(net318),
    .X(_10657_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_427 ();
 sky130_fd_sc_hd__mux4_2 _24824_ (.A0(\w[50][20] ),
    .A1(\w[48][20] ),
    .A2(\w[54][20] ),
    .A3(\w[52][20] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10659_));
 sky130_fd_sc_hd__mux4_2 _24825_ (.A0(\w[58][20] ),
    .A1(\w[56][20] ),
    .A2(\w[62][20] ),
    .A3(\w[60][20] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10660_));
 sky130_fd_sc_hd__mux4_2 _24826_ (.A0(\w[34][20] ),
    .A1(\w[32][20] ),
    .A2(\w[38][20] ),
    .A3(\w[36][20] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10661_));
 sky130_fd_sc_hd__mux4_2 _24827_ (.A0(\w[42][20] ),
    .A1(\w[40][20] ),
    .A2(\w[46][20] ),
    .A3(\w[44][20] ),
    .S0(net372),
    .S1(_00655_),
    .X(_10662_));
 sky130_fd_sc_hd__mux4_2 _24828_ (.A0(_10659_),
    .A1(_10660_),
    .A2(_10661_),
    .A3(_10662_),
    .S0(net325),
    .S1(_10352_),
    .X(_10663_));
 sky130_fd_sc_hd__mux2i_1 _24829_ (.A0(_10657_),
    .A1(_10663_),
    .S(_10373_),
    .Y(_10664_));
 sky130_fd_sc_hd__nand2_1 _24830_ (.A(net348),
    .B(\w[0][20] ),
    .Y(_10665_));
 sky130_fd_sc_hd__o21ai_0 _24831_ (.A1(net287),
    .A2(_10664_),
    .B1(_10665_),
    .Y(_00012_));
 sky130_fd_sc_hd__mux4_2 _24832_ (.A0(\w[18][21] ),
    .A1(\w[16][21] ),
    .A2(\w[22][21] ),
    .A3(\w[20][21] ),
    .S0(net369),
    .S1(net307),
    .X(_10666_));
 sky130_fd_sc_hd__mux4_2 _24833_ (.A0(\w[26][21] ),
    .A1(\w[24][21] ),
    .A2(\w[30][21] ),
    .A3(\w[28][21] ),
    .S0(net369),
    .S1(net307),
    .X(_10667_));
 sky130_fd_sc_hd__mux4_2 _24834_ (.A0(\w[2][21] ),
    .A1(\w[0][21] ),
    .A2(\w[6][21] ),
    .A3(\w[4][21] ),
    .S0(net369),
    .S1(net307),
    .X(_10668_));
 sky130_fd_sc_hd__mux4_2 _24835_ (.A0(\w[10][21] ),
    .A1(\w[8][21] ),
    .A2(\w[14][21] ),
    .A3(\w[12][21] ),
    .S0(net369),
    .S1(net307),
    .X(_10669_));
 sky130_fd_sc_hd__mux4_2 _24836_ (.A0(_10666_),
    .A1(_10667_),
    .A2(_10668_),
    .A3(_10669_),
    .S0(net321),
    .S1(net317),
    .X(_10670_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_426 ();
 sky130_fd_sc_hd__mux4_2 _24838_ (.A0(\w[50][21] ),
    .A1(\w[48][21] ),
    .A2(\w[54][21] ),
    .A3(\w[52][21] ),
    .S0(net370),
    .S1(net306),
    .X(_10672_));
 sky130_fd_sc_hd__mux4_2 _24839_ (.A0(\w[58][21] ),
    .A1(\w[56][21] ),
    .A2(\w[62][21] ),
    .A3(\w[60][21] ),
    .S0(net370),
    .S1(net306),
    .X(_10673_));
 sky130_fd_sc_hd__mux4_2 _24840_ (.A0(\w[34][21] ),
    .A1(\w[32][21] ),
    .A2(\w[38][21] ),
    .A3(\w[36][21] ),
    .S0(net370),
    .S1(net306),
    .X(_10674_));
 sky130_fd_sc_hd__mux4_2 _24841_ (.A0(\w[42][21] ),
    .A1(\w[40][21] ),
    .A2(\w[46][21] ),
    .A3(\w[44][21] ),
    .S0(net370),
    .S1(net306),
    .X(_10675_));
 sky130_fd_sc_hd__mux4_2 _24842_ (.A0(_10672_),
    .A1(_10673_),
    .A2(_10674_),
    .A3(_10675_),
    .S0(net324),
    .S1(net315),
    .X(_10676_));
 sky130_fd_sc_hd__mux2i_1 _24843_ (.A0(_10670_),
    .A1(_10676_),
    .S(net289),
    .Y(_10677_));
 sky130_fd_sc_hd__nand2_1 _24844_ (.A(net348),
    .B(\w[0][21] ),
    .Y(_10678_));
 sky130_fd_sc_hd__o21ai_2 _24845_ (.A1(net286),
    .A2(_10677_),
    .B1(_10678_),
    .Y(_00013_));
 sky130_fd_sc_hd__mux4_2 _24846_ (.A0(\w[18][22] ),
    .A1(\w[16][22] ),
    .A2(\w[22][22] ),
    .A3(\w[20][22] ),
    .S0(net371),
    .S1(net307),
    .X(_10679_));
 sky130_fd_sc_hd__mux4_2 _24847_ (.A0(\w[26][22] ),
    .A1(\w[24][22] ),
    .A2(\w[30][22] ),
    .A3(\w[28][22] ),
    .S0(net371),
    .S1(net307),
    .X(_10680_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_425 ();
 sky130_fd_sc_hd__mux4_2 _24849_ (.A0(\w[2][22] ),
    .A1(\w[0][22] ),
    .A2(\w[6][22] ),
    .A3(\w[4][22] ),
    .S0(net371),
    .S1(net307),
    .X(_10682_));
 sky130_fd_sc_hd__mux4_2 _24850_ (.A0(\w[10][22] ),
    .A1(\w[8][22] ),
    .A2(\w[14][22] ),
    .A3(\w[12][22] ),
    .S0(net371),
    .S1(net307),
    .X(_10683_));
 sky130_fd_sc_hd__mux4_2 _24851_ (.A0(_10679_),
    .A1(_10680_),
    .A2(_10682_),
    .A3(_10683_),
    .S0(net320),
    .S1(net316),
    .X(_10684_));
 sky130_fd_sc_hd__mux4_2 _24852_ (.A0(\w[50][22] ),
    .A1(\w[48][22] ),
    .A2(\w[54][22] ),
    .A3(\w[52][22] ),
    .S0(net372),
    .S1(net303),
    .X(_10685_));
 sky130_fd_sc_hd__mux4_2 _24853_ (.A0(\w[58][22] ),
    .A1(\w[56][22] ),
    .A2(\w[62][22] ),
    .A3(\w[60][22] ),
    .S0(net372),
    .S1(net303),
    .X(_10686_));
 sky130_fd_sc_hd__mux4_2 _24854_ (.A0(\w[34][22] ),
    .A1(\w[32][22] ),
    .A2(\w[38][22] ),
    .A3(\w[36][22] ),
    .S0(net372),
    .S1(net303),
    .X(_10687_));
 sky130_fd_sc_hd__mux4_2 _24855_ (.A0(\w[42][22] ),
    .A1(\w[40][22] ),
    .A2(\w[46][22] ),
    .A3(\w[44][22] ),
    .S0(net372),
    .S1(net303),
    .X(_10688_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_424 ();
 sky130_fd_sc_hd__mux4_2 _24857_ (.A0(_10685_),
    .A1(_10686_),
    .A2(_10687_),
    .A3(_10688_),
    .S0(net321),
    .S1(net317),
    .X(_10690_));
 sky130_fd_sc_hd__mux2i_1 _24858_ (.A0(_10684_),
    .A1(_10690_),
    .S(net289),
    .Y(_10691_));
 sky130_fd_sc_hd__nand2_1 _24859_ (.A(net348),
    .B(\w[0][22] ),
    .Y(_10692_));
 sky130_fd_sc_hd__o21ai_2 _24860_ (.A1(net287),
    .A2(_10691_),
    .B1(_10692_),
    .Y(_00014_));
 sky130_fd_sc_hd__mux4_2 _24861_ (.A0(\w[18][23] ),
    .A1(\w[16][23] ),
    .A2(\w[22][23] ),
    .A3(\w[20][23] ),
    .S0(net367),
    .S1(net303),
    .X(_10693_));
 sky130_fd_sc_hd__mux4_2 _24862_ (.A0(\w[26][23] ),
    .A1(\w[24][23] ),
    .A2(\w[30][23] ),
    .A3(\w[28][23] ),
    .S0(net367),
    .S1(net303),
    .X(_10694_));
 sky130_fd_sc_hd__mux4_2 _24863_ (.A0(\w[2][23] ),
    .A1(\w[0][23] ),
    .A2(\w[6][23] ),
    .A3(\w[4][23] ),
    .S0(net367),
    .S1(net305),
    .X(_10695_));
 sky130_fd_sc_hd__mux4_2 _24864_ (.A0(\w[10][23] ),
    .A1(\w[8][23] ),
    .A2(\w[14][23] ),
    .A3(\w[12][23] ),
    .S0(net367),
    .S1(net303),
    .X(_10696_));
 sky130_fd_sc_hd__mux4_2 _24865_ (.A0(_10693_),
    .A1(_10694_),
    .A2(_10695_),
    .A3(_10696_),
    .S0(net322),
    .S1(net313),
    .X(_10697_));
 sky130_fd_sc_hd__mux4_2 _24866_ (.A0(\w[50][23] ),
    .A1(\w[48][23] ),
    .A2(\w[54][23] ),
    .A3(\w[52][23] ),
    .S0(net366),
    .S1(net306),
    .X(_10698_));
 sky130_fd_sc_hd__mux4_2 _24867_ (.A0(\w[58][23] ),
    .A1(\w[56][23] ),
    .A2(\w[62][23] ),
    .A3(\w[60][23] ),
    .S0(net366),
    .S1(net306),
    .X(_10699_));
 sky130_fd_sc_hd__mux4_2 _24868_ (.A0(\w[34][23] ),
    .A1(\w[32][23] ),
    .A2(\w[38][23] ),
    .A3(\w[36][23] ),
    .S0(net366),
    .S1(net306),
    .X(_10700_));
 sky130_fd_sc_hd__mux4_2 _24869_ (.A0(\w[42][23] ),
    .A1(\w[40][23] ),
    .A2(\w[46][23] ),
    .A3(\w[44][23] ),
    .S0(net366),
    .S1(net306),
    .X(_10701_));
 sky130_fd_sc_hd__mux4_2 _24870_ (.A0(_10698_),
    .A1(_10699_),
    .A2(_10700_),
    .A3(_10701_),
    .S0(net324),
    .S1(net313),
    .X(_10702_));
 sky130_fd_sc_hd__mux2i_1 _24871_ (.A0(_10697_),
    .A1(_10702_),
    .S(net288),
    .Y(_10703_));
 sky130_fd_sc_hd__nand2_1 _24872_ (.A(net348),
    .B(\w[0][23] ),
    .Y(_10704_));
 sky130_fd_sc_hd__o21ai_1 _24873_ (.A1(net286),
    .A2(_10703_),
    .B1(_10704_),
    .Y(_00015_));
 sky130_fd_sc_hd__mux4_2 _24874_ (.A0(\w[18][24] ),
    .A1(\w[16][24] ),
    .A2(\w[22][24] ),
    .A3(\w[20][24] ),
    .S0(net371),
    .S1(net307),
    .X(_10705_));
 sky130_fd_sc_hd__mux4_2 _24875_ (.A0(\w[26][24] ),
    .A1(\w[24][24] ),
    .A2(\w[30][24] ),
    .A3(\w[28][24] ),
    .S0(net371),
    .S1(net307),
    .X(_10706_));
 sky130_fd_sc_hd__mux4_2 _24876_ (.A0(\w[2][24] ),
    .A1(\w[0][24] ),
    .A2(\w[6][24] ),
    .A3(\w[4][24] ),
    .S0(net371),
    .S1(net307),
    .X(_10707_));
 sky130_fd_sc_hd__mux4_2 _24877_ (.A0(\w[10][24] ),
    .A1(\w[8][24] ),
    .A2(\w[14][24] ),
    .A3(\w[12][24] ),
    .S0(net371),
    .S1(net307),
    .X(_10708_));
 sky130_fd_sc_hd__mux4_2 _24878_ (.A0(_10705_),
    .A1(_10706_),
    .A2(_10707_),
    .A3(_10708_),
    .S0(net320),
    .S1(net316),
    .X(_10709_));
 sky130_fd_sc_hd__mux4_2 _24879_ (.A0(\w[50][24] ),
    .A1(\w[48][24] ),
    .A2(\w[54][24] ),
    .A3(\w[52][24] ),
    .S0(net369),
    .S1(net303),
    .X(_10710_));
 sky130_fd_sc_hd__mux4_2 _24880_ (.A0(\w[58][24] ),
    .A1(\w[56][24] ),
    .A2(\w[62][24] ),
    .A3(\w[60][24] ),
    .S0(net369),
    .S1(net303),
    .X(_10711_));
 sky130_fd_sc_hd__mux4_2 _24881_ (.A0(\w[34][24] ),
    .A1(\w[32][24] ),
    .A2(\w[38][24] ),
    .A3(\w[36][24] ),
    .S0(net369),
    .S1(net303),
    .X(_10712_));
 sky130_fd_sc_hd__mux4_2 _24882_ (.A0(\w[42][24] ),
    .A1(\w[40][24] ),
    .A2(\w[46][24] ),
    .A3(\w[44][24] ),
    .S0(net369),
    .S1(net303),
    .X(_10713_));
 sky130_fd_sc_hd__mux4_2 _24883_ (.A0(_10710_),
    .A1(_10711_),
    .A2(_10712_),
    .A3(_10713_),
    .S0(net321),
    .S1(net317),
    .X(_10714_));
 sky130_fd_sc_hd__mux2i_1 _24884_ (.A0(_10709_),
    .A1(_10714_),
    .S(net290),
    .Y(_10715_));
 sky130_fd_sc_hd__nand2_1 _24885_ (.A(net348),
    .B(\w[0][24] ),
    .Y(_10716_));
 sky130_fd_sc_hd__o21ai_2 _24886_ (.A1(net287),
    .A2(_10715_),
    .B1(_10716_),
    .Y(_00016_));
 sky130_fd_sc_hd__mux4_2 _24887_ (.A0(\w[18][25] ),
    .A1(\w[16][25] ),
    .A2(\w[22][25] ),
    .A3(\w[20][25] ),
    .S0(net369),
    .S1(net303),
    .X(_10717_));
 sky130_fd_sc_hd__mux4_2 _24888_ (.A0(\w[26][25] ),
    .A1(\w[24][25] ),
    .A2(\w[30][25] ),
    .A3(\w[28][25] ),
    .S0(net369),
    .S1(net303),
    .X(_10718_));
 sky130_fd_sc_hd__mux4_2 _24889_ (.A0(\w[2][25] ),
    .A1(\w[0][25] ),
    .A2(\w[6][25] ),
    .A3(\w[4][25] ),
    .S0(net369),
    .S1(net303),
    .X(_10719_));
 sky130_fd_sc_hd__mux4_2 _24890_ (.A0(\w[10][25] ),
    .A1(\w[8][25] ),
    .A2(\w[14][25] ),
    .A3(\w[12][25] ),
    .S0(net369),
    .S1(net303),
    .X(_10720_));
 sky130_fd_sc_hd__mux4_2 _24891_ (.A0(_10717_),
    .A1(_10718_),
    .A2(_10719_),
    .A3(_10720_),
    .S0(net321),
    .S1(net317),
    .X(_10721_));
 sky130_fd_sc_hd__mux4_2 _24892_ (.A0(\w[50][25] ),
    .A1(\w[48][25] ),
    .A2(\w[54][25] ),
    .A3(\w[52][25] ),
    .S0(net368),
    .S1(net305),
    .X(_10722_));
 sky130_fd_sc_hd__mux4_2 _24893_ (.A0(\w[58][25] ),
    .A1(\w[56][25] ),
    .A2(\w[62][25] ),
    .A3(\w[60][25] ),
    .S0(net368),
    .S1(net305),
    .X(_10723_));
 sky130_fd_sc_hd__mux4_2 _24894_ (.A0(\w[34][25] ),
    .A1(\w[32][25] ),
    .A2(\w[38][25] ),
    .A3(\w[36][25] ),
    .S0(net368),
    .S1(net305),
    .X(_10724_));
 sky130_fd_sc_hd__mux4_2 _24895_ (.A0(\w[42][25] ),
    .A1(\w[40][25] ),
    .A2(\w[46][25] ),
    .A3(\w[44][25] ),
    .S0(net368),
    .S1(net305),
    .X(_10725_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_423 ();
 sky130_fd_sc_hd__mux4_2 _24897_ (.A0(_10722_),
    .A1(_10723_),
    .A2(_10724_),
    .A3(_10725_),
    .S0(net324),
    .S1(net315),
    .X(_10727_));
 sky130_fd_sc_hd__mux2i_1 _24898_ (.A0(_10721_),
    .A1(_10727_),
    .S(net289),
    .Y(_10728_));
 sky130_fd_sc_hd__nand2_2 _24899_ (.A(net348),
    .B(\w[0][25] ),
    .Y(_10729_));
 sky130_fd_sc_hd__o21ai_4 _24900_ (.A1(net286),
    .A2(_10728_),
    .B1(_10729_),
    .Y(_00017_));
 sky130_fd_sc_hd__mux4_2 _24901_ (.A0(\w[18][26] ),
    .A1(\w[16][26] ),
    .A2(\w[22][26] ),
    .A3(\w[20][26] ),
    .S0(net369),
    .S1(net307),
    .X(_10730_));
 sky130_fd_sc_hd__mux4_2 _24902_ (.A0(\w[26][26] ),
    .A1(\w[24][26] ),
    .A2(\w[30][26] ),
    .A3(\w[28][26] ),
    .S0(net369),
    .S1(net307),
    .X(_10731_));
 sky130_fd_sc_hd__mux4_2 _24903_ (.A0(\w[2][26] ),
    .A1(\w[0][26] ),
    .A2(\w[6][26] ),
    .A3(\w[4][26] ),
    .S0(net369),
    .S1(net307),
    .X(_10732_));
 sky130_fd_sc_hd__mux4_2 _24904_ (.A0(\w[10][26] ),
    .A1(\w[8][26] ),
    .A2(\w[14][26] ),
    .A3(\w[12][26] ),
    .S0(net369),
    .S1(net307),
    .X(_10733_));
 sky130_fd_sc_hd__mux4_2 _24905_ (.A0(_10730_),
    .A1(_10731_),
    .A2(_10732_),
    .A3(_10733_),
    .S0(net321),
    .S1(net317),
    .X(_10734_));
 sky130_fd_sc_hd__mux4_2 _24906_ (.A0(\w[50][26] ),
    .A1(\w[48][26] ),
    .A2(\w[54][26] ),
    .A3(\w[52][26] ),
    .S0(net369),
    .S1(net303),
    .X(_10735_));
 sky130_fd_sc_hd__mux4_2 _24907_ (.A0(\w[58][26] ),
    .A1(\w[56][26] ),
    .A2(\w[62][26] ),
    .A3(\w[60][26] ),
    .S0(net369),
    .S1(net303),
    .X(_10736_));
 sky130_fd_sc_hd__mux4_2 _24908_ (.A0(\w[34][26] ),
    .A1(\w[32][26] ),
    .A2(\w[38][26] ),
    .A3(\w[36][26] ),
    .S0(net369),
    .S1(net303),
    .X(_10737_));
 sky130_fd_sc_hd__mux4_2 _24909_ (.A0(\w[42][26] ),
    .A1(\w[40][26] ),
    .A2(\w[46][26] ),
    .A3(\w[44][26] ),
    .S0(net369),
    .S1(net303),
    .X(_10738_));
 sky130_fd_sc_hd__mux4_2 _24910_ (.A0(_10735_),
    .A1(_10736_),
    .A2(_10737_),
    .A3(_10738_),
    .S0(net321),
    .S1(net317),
    .X(_10739_));
 sky130_fd_sc_hd__mux2i_1 _24911_ (.A0(_10734_),
    .A1(_10739_),
    .S(net289),
    .Y(_10740_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_422 ();
 sky130_fd_sc_hd__nand2_2 _24913_ (.A(net348),
    .B(\w[0][26] ),
    .Y(_10742_));
 sky130_fd_sc_hd__o21ai_4 _24914_ (.A1(net286),
    .A2(_10740_),
    .B1(_10742_),
    .Y(_00018_));
 sky130_fd_sc_hd__mux4_2 _24915_ (.A0(\w[18][27] ),
    .A1(\w[16][27] ),
    .A2(\w[22][27] ),
    .A3(\w[20][27] ),
    .S0(net367),
    .S1(net303),
    .X(_10743_));
 sky130_fd_sc_hd__mux4_2 _24916_ (.A0(\w[26][27] ),
    .A1(\w[24][27] ),
    .A2(\w[30][27] ),
    .A3(\w[28][27] ),
    .S0(net367),
    .S1(net303),
    .X(_10744_));
 sky130_fd_sc_hd__mux4_2 _24917_ (.A0(\w[2][27] ),
    .A1(\w[0][27] ),
    .A2(\w[6][27] ),
    .A3(\w[4][27] ),
    .S0(net367),
    .S1(net303),
    .X(_10745_));
 sky130_fd_sc_hd__mux4_2 _24918_ (.A0(\w[10][27] ),
    .A1(\w[8][27] ),
    .A2(\w[14][27] ),
    .A3(\w[12][27] ),
    .S0(net367),
    .S1(net303),
    .X(_10746_));
 sky130_fd_sc_hd__mux4_2 _24919_ (.A0(_10743_),
    .A1(_10744_),
    .A2(_10745_),
    .A3(_10746_),
    .S0(net322),
    .S1(net313),
    .X(_10747_));
 sky130_fd_sc_hd__mux4_2 _24920_ (.A0(\w[50][27] ),
    .A1(\w[48][27] ),
    .A2(\w[54][27] ),
    .A3(\w[52][27] ),
    .S0(net368),
    .S1(net305),
    .X(_10748_));
 sky130_fd_sc_hd__mux4_2 _24921_ (.A0(\w[58][27] ),
    .A1(\w[56][27] ),
    .A2(\w[62][27] ),
    .A3(\w[60][27] ),
    .S0(net368),
    .S1(net305),
    .X(_10749_));
 sky130_fd_sc_hd__mux4_2 _24922_ (.A0(\w[34][27] ),
    .A1(\w[32][27] ),
    .A2(\w[38][27] ),
    .A3(\w[36][27] ),
    .S0(net368),
    .S1(net305),
    .X(_10750_));
 sky130_fd_sc_hd__mux4_2 _24923_ (.A0(\w[42][27] ),
    .A1(\w[40][27] ),
    .A2(\w[46][27] ),
    .A3(\w[44][27] ),
    .S0(net368),
    .S1(net305),
    .X(_10751_));
 sky130_fd_sc_hd__mux4_2 _24924_ (.A0(_10748_),
    .A1(_10749_),
    .A2(_10750_),
    .A3(_10751_),
    .S0(net322),
    .S1(net313),
    .X(_10752_));
 sky130_fd_sc_hd__mux2i_1 _24925_ (.A0(_10747_),
    .A1(_10752_),
    .S(net288),
    .Y(_10753_));
 sky130_fd_sc_hd__nand2_2 _24926_ (.A(net348),
    .B(\w[0][27] ),
    .Y(_10754_));
 sky130_fd_sc_hd__o21ai_4 _24927_ (.A1(net286),
    .A2(_10753_),
    .B1(_10754_),
    .Y(_00019_));
 sky130_fd_sc_hd__mux4_2 _24928_ (.A0(\w[18][28] ),
    .A1(\w[16][28] ),
    .A2(\w[22][28] ),
    .A3(\w[20][28] ),
    .S0(net367),
    .S1(net303),
    .X(_10755_));
 sky130_fd_sc_hd__mux4_2 _24929_ (.A0(\w[26][28] ),
    .A1(\w[24][28] ),
    .A2(\w[30][28] ),
    .A3(\w[28][28] ),
    .S0(net367),
    .S1(net303),
    .X(_10756_));
 sky130_fd_sc_hd__mux4_2 _24930_ (.A0(\w[2][28] ),
    .A1(\w[0][28] ),
    .A2(\w[6][28] ),
    .A3(\w[4][28] ),
    .S0(net367),
    .S1(net303),
    .X(_10757_));
 sky130_fd_sc_hd__mux4_2 _24931_ (.A0(\w[10][28] ),
    .A1(\w[8][28] ),
    .A2(\w[14][28] ),
    .A3(\w[12][28] ),
    .S0(net367),
    .S1(net303),
    .X(_10758_));
 sky130_fd_sc_hd__mux4_2 _24932_ (.A0(_10755_),
    .A1(_10756_),
    .A2(_10757_),
    .A3(_10758_),
    .S0(net322),
    .S1(net313),
    .X(_10759_));
 sky130_fd_sc_hd__mux4_2 _24933_ (.A0(\w[50][28] ),
    .A1(\w[48][28] ),
    .A2(\w[54][28] ),
    .A3(\w[52][28] ),
    .S0(net368),
    .S1(net305),
    .X(_10760_));
 sky130_fd_sc_hd__mux4_2 _24934_ (.A0(\w[58][28] ),
    .A1(\w[56][28] ),
    .A2(\w[62][28] ),
    .A3(\w[60][28] ),
    .S0(net368),
    .S1(net305),
    .X(_10761_));
 sky130_fd_sc_hd__mux4_2 _24935_ (.A0(\w[34][28] ),
    .A1(\w[32][28] ),
    .A2(\w[38][28] ),
    .A3(\w[36][28] ),
    .S0(net368),
    .S1(net305),
    .X(_10762_));
 sky130_fd_sc_hd__mux4_2 _24936_ (.A0(\w[42][28] ),
    .A1(\w[40][28] ),
    .A2(\w[46][28] ),
    .A3(\w[44][28] ),
    .S0(net368),
    .S1(net305),
    .X(_10763_));
 sky130_fd_sc_hd__mux4_2 _24937_ (.A0(_10760_),
    .A1(_10761_),
    .A2(_10762_),
    .A3(_10763_),
    .S0(net322),
    .S1(net313),
    .X(_10764_));
 sky130_fd_sc_hd__mux2i_1 _24938_ (.A0(_10759_),
    .A1(_10764_),
    .S(net288),
    .Y(_10765_));
 sky130_fd_sc_hd__nand2_2 _24939_ (.A(net348),
    .B(\w[0][28] ),
    .Y(_10766_));
 sky130_fd_sc_hd__o21ai_4 _24940_ (.A1(net286),
    .A2(_10765_),
    .B1(_10766_),
    .Y(_00020_));
 sky130_fd_sc_hd__mux4_2 _24941_ (.A0(\w[18][29] ),
    .A1(\w[16][29] ),
    .A2(\w[22][29] ),
    .A3(\w[20][29] ),
    .S0(net367),
    .S1(net303),
    .X(_10767_));
 sky130_fd_sc_hd__mux4_2 _24942_ (.A0(\w[26][29] ),
    .A1(\w[24][29] ),
    .A2(\w[30][29] ),
    .A3(\w[28][29] ),
    .S0(net367),
    .S1(net303),
    .X(_10768_));
 sky130_fd_sc_hd__mux4_2 _24943_ (.A0(\w[2][29] ),
    .A1(\w[0][29] ),
    .A2(\w[6][29] ),
    .A3(\w[4][29] ),
    .S0(net367),
    .S1(net303),
    .X(_10769_));
 sky130_fd_sc_hd__mux4_2 _24944_ (.A0(\w[10][29] ),
    .A1(\w[8][29] ),
    .A2(\w[14][29] ),
    .A3(\w[12][29] ),
    .S0(net367),
    .S1(net303),
    .X(_10770_));
 sky130_fd_sc_hd__mux4_2 _24945_ (.A0(_10767_),
    .A1(_10768_),
    .A2(_10769_),
    .A3(_10770_),
    .S0(net322),
    .S1(net313),
    .X(_10771_));
 sky130_fd_sc_hd__mux4_2 _24946_ (.A0(\w[50][29] ),
    .A1(\w[48][29] ),
    .A2(\w[54][29] ),
    .A3(\w[52][29] ),
    .S0(net368),
    .S1(net305),
    .X(_10772_));
 sky130_fd_sc_hd__mux4_2 _24947_ (.A0(\w[58][29] ),
    .A1(\w[56][29] ),
    .A2(\w[62][29] ),
    .A3(\w[60][29] ),
    .S0(net368),
    .S1(net305),
    .X(_10773_));
 sky130_fd_sc_hd__mux4_2 _24948_ (.A0(\w[34][29] ),
    .A1(\w[32][29] ),
    .A2(\w[38][29] ),
    .A3(\w[36][29] ),
    .S0(net368),
    .S1(net305),
    .X(_10774_));
 sky130_fd_sc_hd__mux4_2 _24949_ (.A0(\w[42][29] ),
    .A1(\w[40][29] ),
    .A2(\w[46][29] ),
    .A3(\w[44][29] ),
    .S0(net368),
    .S1(net305),
    .X(_10775_));
 sky130_fd_sc_hd__mux4_2 _24950_ (.A0(_10772_),
    .A1(_10773_),
    .A2(_10774_),
    .A3(_10775_),
    .S0(net322),
    .S1(net313),
    .X(_10776_));
 sky130_fd_sc_hd__mux2i_1 _24951_ (.A0(_10771_),
    .A1(_10776_),
    .S(net288),
    .Y(_10777_));
 sky130_fd_sc_hd__nand2_2 _24952_ (.A(reset_hash),
    .B(\w[0][29] ),
    .Y(_10778_));
 sky130_fd_sc_hd__o21ai_4 _24953_ (.A1(net286),
    .A2(_10777_),
    .B1(_10778_),
    .Y(_00021_));
 sky130_fd_sc_hd__mux4_2 _24954_ (.A0(\w[18][30] ),
    .A1(\w[16][30] ),
    .A2(\w[22][30] ),
    .A3(\w[20][30] ),
    .S0(net367),
    .S1(net303),
    .X(_10779_));
 sky130_fd_sc_hd__mux4_2 _24955_ (.A0(\w[26][30] ),
    .A1(\w[24][30] ),
    .A2(\w[30][30] ),
    .A3(\w[28][30] ),
    .S0(net367),
    .S1(net303),
    .X(_10780_));
 sky130_fd_sc_hd__mux4_2 _24956_ (.A0(\w[2][30] ),
    .A1(\w[0][30] ),
    .A2(\w[6][30] ),
    .A3(\w[4][30] ),
    .S0(net367),
    .S1(net303),
    .X(_10781_));
 sky130_fd_sc_hd__mux4_2 _24957_ (.A0(\w[10][30] ),
    .A1(\w[8][30] ),
    .A2(\w[14][30] ),
    .A3(\w[12][30] ),
    .S0(net367),
    .S1(net303),
    .X(_10782_));
 sky130_fd_sc_hd__mux4_2 _24958_ (.A0(_10779_),
    .A1(_10780_),
    .A2(_10781_),
    .A3(_10782_),
    .S0(net322),
    .S1(net313),
    .X(_10783_));
 sky130_fd_sc_hd__mux4_2 _24959_ (.A0(\w[50][30] ),
    .A1(\w[48][30] ),
    .A2(\w[54][30] ),
    .A3(\w[52][30] ),
    .S0(net368),
    .S1(net305),
    .X(_10784_));
 sky130_fd_sc_hd__mux4_2 _24960_ (.A0(\w[58][30] ),
    .A1(\w[56][30] ),
    .A2(\w[62][30] ),
    .A3(\w[60][30] ),
    .S0(net368),
    .S1(net305),
    .X(_10785_));
 sky130_fd_sc_hd__mux4_2 _24961_ (.A0(\w[34][30] ),
    .A1(\w[32][30] ),
    .A2(\w[38][30] ),
    .A3(\w[36][30] ),
    .S0(net368),
    .S1(net305),
    .X(_10786_));
 sky130_fd_sc_hd__mux4_2 _24962_ (.A0(\w[42][30] ),
    .A1(\w[40][30] ),
    .A2(\w[46][30] ),
    .A3(\w[44][30] ),
    .S0(net368),
    .S1(net305),
    .X(_10787_));
 sky130_fd_sc_hd__mux4_2 _24963_ (.A0(_10784_),
    .A1(_10785_),
    .A2(_10786_),
    .A3(_10787_),
    .S0(net322),
    .S1(net313),
    .X(_10788_));
 sky130_fd_sc_hd__mux2i_1 _24964_ (.A0(_10783_),
    .A1(_10788_),
    .S(net288),
    .Y(_10789_));
 sky130_fd_sc_hd__nand2_2 _24965_ (.A(reset_hash),
    .B(\w[0][30] ),
    .Y(_10790_));
 sky130_fd_sc_hd__o21ai_4 _24966_ (.A1(net286),
    .A2(_10789_),
    .B1(_10790_),
    .Y(_00023_));
 sky130_fd_sc_hd__mux4_2 _24967_ (.A0(\w[18][31] ),
    .A1(\w[16][31] ),
    .A2(\w[22][31] ),
    .A3(\w[20][31] ),
    .S0(net369),
    .S1(net303),
    .X(_10791_));
 sky130_fd_sc_hd__mux4_2 _24968_ (.A0(\w[26][31] ),
    .A1(\w[24][31] ),
    .A2(\w[30][31] ),
    .A3(\w[28][31] ),
    .S0(net369),
    .S1(net303),
    .X(_10792_));
 sky130_fd_sc_hd__mux4_2 _24969_ (.A0(\w[2][31] ),
    .A1(\w[0][31] ),
    .A2(\w[6][31] ),
    .A3(\w[4][31] ),
    .S0(net369),
    .S1(net303),
    .X(_10793_));
 sky130_fd_sc_hd__mux4_2 _24970_ (.A0(\w[10][31] ),
    .A1(\w[8][31] ),
    .A2(\w[14][31] ),
    .A3(\w[12][31] ),
    .S0(net369),
    .S1(net303),
    .X(_10794_));
 sky130_fd_sc_hd__mux4_2 _24971_ (.A0(_10791_),
    .A1(_10792_),
    .A2(_10793_),
    .A3(_10794_),
    .S0(net321),
    .S1(net317),
    .X(_10795_));
 sky130_fd_sc_hd__mux4_2 _24972_ (.A0(\w[50][31] ),
    .A1(\w[48][31] ),
    .A2(\w[54][31] ),
    .A3(\w[52][31] ),
    .S0(net370),
    .S1(net306),
    .X(_10796_));
 sky130_fd_sc_hd__mux4_2 _24973_ (.A0(\w[58][31] ),
    .A1(\w[56][31] ),
    .A2(\w[62][31] ),
    .A3(\w[60][31] ),
    .S0(net370),
    .S1(net306),
    .X(_10797_));
 sky130_fd_sc_hd__mux4_2 _24974_ (.A0(\w[34][31] ),
    .A1(\w[32][31] ),
    .A2(\w[38][31] ),
    .A3(\w[36][31] ),
    .S0(net370),
    .S1(net306),
    .X(_10798_));
 sky130_fd_sc_hd__mux4_2 _24975_ (.A0(\w[42][31] ),
    .A1(\w[40][31] ),
    .A2(\w[46][31] ),
    .A3(\w[44][31] ),
    .S0(net370),
    .S1(net306),
    .X(_10799_));
 sky130_fd_sc_hd__mux4_2 _24976_ (.A0(_10796_),
    .A1(_10797_),
    .A2(_10798_),
    .A3(_10799_),
    .S0(net324),
    .S1(net315),
    .X(_10800_));
 sky130_fd_sc_hd__mux2i_1 _24977_ (.A0(_10795_),
    .A1(_10800_),
    .S(net289),
    .Y(_10801_));
 sky130_fd_sc_hd__nand2_2 _24978_ (.A(net348),
    .B(\w[0][31] ),
    .Y(_10802_));
 sky130_fd_sc_hd__o21ai_4 _24979_ (.A1(net286),
    .A2(_10801_),
    .B1(_10802_),
    .Y(_00024_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_413 ();
 sky130_fd_sc_hd__mux4_2 _24989_ (.A0(\w[1][3] ),
    .A1(\w[5][3] ),
    .A2(\w[3][3] ),
    .A3(\w[7][3] ),
    .S0(net519),
    .S1(net528),
    .X(_10812_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_409 ();
 sky130_fd_sc_hd__mux4_2 _24994_ (.A0(\w[9][3] ),
    .A1(\w[13][3] ),
    .A2(\w[11][3] ),
    .A3(\w[15][3] ),
    .S0(net519),
    .S1(net528),
    .X(_10817_));
 sky130_fd_sc_hd__mux4_2 _24995_ (.A0(\w[17][3] ),
    .A1(\w[21][3] ),
    .A2(\w[19][3] ),
    .A3(\w[23][3] ),
    .S0(net519),
    .S1(net528),
    .X(_10818_));
 sky130_fd_sc_hd__mux4_2 _24996_ (.A0(\w[25][3] ),
    .A1(\w[29][3] ),
    .A2(\w[27][3] ),
    .A3(\w[31][3] ),
    .S0(net519),
    .S1(net528),
    .X(_10819_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_404 ();
 sky130_fd_sc_hd__mux4_2 _25002_ (.A0(_10812_),
    .A1(_10817_),
    .A2(_10818_),
    .A3(_10819_),
    .S0(net518),
    .S1(net549),
    .X(_10825_));
 sky130_fd_sc_hd__mux4_2 _25003_ (.A0(\w[33][3] ),
    .A1(\w[37][3] ),
    .A2(\w[35][3] ),
    .A3(\w[39][3] ),
    .S0(net519),
    .S1(net528),
    .X(_10826_));
 sky130_fd_sc_hd__mux4_2 _25004_ (.A0(\w[41][3] ),
    .A1(\w[45][3] ),
    .A2(\w[43][3] ),
    .A3(\w[47][3] ),
    .S0(net519),
    .S1(net528),
    .X(_10827_));
 sky130_fd_sc_hd__mux4_2 _25005_ (.A0(\w[49][3] ),
    .A1(\w[53][3] ),
    .A2(\w[51][3] ),
    .A3(\w[55][3] ),
    .S0(net519),
    .S1(net528),
    .X(_10828_));
 sky130_fd_sc_hd__mux4_2 _25006_ (.A0(\w[57][3] ),
    .A1(\w[61][3] ),
    .A2(\w[59][3] ),
    .A3(\w[63][3] ),
    .S0(net519),
    .S1(net528),
    .X(_10829_));
 sky130_fd_sc_hd__mux4_2 _25007_ (.A0(_10826_),
    .A1(_10827_),
    .A2(_10828_),
    .A3(_10829_),
    .S0(net518),
    .S1(net549),
    .X(_10830_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_402 ();
 sky130_fd_sc_hd__mux2i_4 _25010_ (.A0(_10825_),
    .A1(_10830_),
    .S(net513),
    .Y(_10833_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_399 ();
 sky130_fd_sc_hd__mux4_2 _25014_ (.A0(\w[1][18] ),
    .A1(\w[5][18] ),
    .A2(\w[3][18] ),
    .A3(\w[7][18] ),
    .S0(net524),
    .S1(net529),
    .X(_10837_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_397 ();
 sky130_fd_sc_hd__mux4_2 _25017_ (.A0(\w[9][18] ),
    .A1(\w[13][18] ),
    .A2(\w[11][18] ),
    .A3(\w[15][18] ),
    .S0(net524),
    .S1(net529),
    .X(_10840_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_395 ();
 sky130_fd_sc_hd__mux4_2 _25020_ (.A0(\w[17][18] ),
    .A1(\w[21][18] ),
    .A2(\w[19][18] ),
    .A3(\w[23][18] ),
    .S0(net524),
    .S1(net529),
    .X(_10843_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_393 ();
 sky130_fd_sc_hd__mux4_2 _25023_ (.A0(\w[25][18] ),
    .A1(\w[29][18] ),
    .A2(\w[27][18] ),
    .A3(\w[31][18] ),
    .S0(net524),
    .S1(net529),
    .X(_10846_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_391 ();
 sky130_fd_sc_hd__mux4_2 _25026_ (.A0(_10837_),
    .A1(_10840_),
    .A2(_10843_),
    .A3(_10846_),
    .S0(net517),
    .S1(net515),
    .X(_10849_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_390 ();
 sky130_fd_sc_hd__mux4_2 _25028_ (.A0(\w[33][18] ),
    .A1(\w[37][18] ),
    .A2(\w[35][18] ),
    .A3(\w[39][18] ),
    .S0(net524),
    .S1(net530),
    .X(_10851_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_388 ();
 sky130_fd_sc_hd__mux4_2 _25031_ (.A0(\w[41][18] ),
    .A1(\w[45][18] ),
    .A2(\w[43][18] ),
    .A3(\w[47][18] ),
    .S0(net525),
    .S1(net530),
    .X(_10854_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_386 ();
 sky130_fd_sc_hd__mux4_2 _25034_ (.A0(\w[49][18] ),
    .A1(\w[53][18] ),
    .A2(\w[51][18] ),
    .A3(\w[55][18] ),
    .S0(net525),
    .S1(net530),
    .X(_10857_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_384 ();
 sky130_fd_sc_hd__mux4_2 _25037_ (.A0(\w[57][18] ),
    .A1(\w[61][18] ),
    .A2(\w[59][18] ),
    .A3(\w[63][18] ),
    .S0(net525),
    .S1(net530),
    .X(_10860_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_382 ();
 sky130_fd_sc_hd__mux4_2 _25040_ (.A0(_10851_),
    .A1(_10854_),
    .A2(_10857_),
    .A3(_10860_),
    .S0(net517),
    .S1(net515),
    .X(_10863_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_381 ();
 sky130_fd_sc_hd__mux2i_4 _25042_ (.A0(_10849_),
    .A1(_10863_),
    .S(\count15_1[5] ),
    .Y(_10865_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_379 ();
 sky130_fd_sc_hd__mux4_2 _25045_ (.A0(\w[1][7] ),
    .A1(\w[5][7] ),
    .A2(\w[3][7] ),
    .A3(\w[7][7] ),
    .S0(net519),
    .S1(net532),
    .X(_10868_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_377 ();
 sky130_fd_sc_hd__mux4_2 _25048_ (.A0(\w[9][7] ),
    .A1(\w[13][7] ),
    .A2(\w[11][7] ),
    .A3(\w[15][7] ),
    .S0(net519),
    .S1(net532),
    .X(_10871_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_376 ();
 sky130_fd_sc_hd__mux4_2 _25050_ (.A0(\w[17][7] ),
    .A1(\w[21][7] ),
    .A2(\w[19][7] ),
    .A3(\w[23][7] ),
    .S0(net519),
    .S1(net532),
    .X(_10873_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_375 ();
 sky130_fd_sc_hd__mux4_2 _25052_ (.A0(\w[25][7] ),
    .A1(\w[29][7] ),
    .A2(\w[27][7] ),
    .A3(\w[31][7] ),
    .S0(net519),
    .S1(net532),
    .X(_10875_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_373 ();
 sky130_fd_sc_hd__mux4_2 _25055_ (.A0(_10868_),
    .A1(_10871_),
    .A2(_10873_),
    .A3(_10875_),
    .S0(net518),
    .S1(net549),
    .X(_10878_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_371 ();
 sky130_fd_sc_hd__mux4_2 _25058_ (.A0(\w[33][7] ),
    .A1(\w[37][7] ),
    .A2(\w[35][7] ),
    .A3(\w[39][7] ),
    .S0(net519),
    .S1(net531),
    .X(_10881_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_369 ();
 sky130_fd_sc_hd__mux4_2 _25061_ (.A0(\w[41][7] ),
    .A1(\w[45][7] ),
    .A2(\w[43][7] ),
    .A3(\w[47][7] ),
    .S0(net519),
    .S1(net531),
    .X(_10884_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_368 ();
 sky130_fd_sc_hd__mux4_2 _25063_ (.A0(\w[49][7] ),
    .A1(\w[53][7] ),
    .A2(\w[51][7] ),
    .A3(\w[55][7] ),
    .S0(net519),
    .S1(net531),
    .X(_10886_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_366 ();
 sky130_fd_sc_hd__mux4_2 _25066_ (.A0(\w[57][7] ),
    .A1(\w[61][7] ),
    .A2(\w[59][7] ),
    .A3(\w[63][7] ),
    .S0(net519),
    .S1(net531),
    .X(_10889_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_364 ();
 sky130_fd_sc_hd__mux4_2 _25069_ (.A0(_10881_),
    .A1(_10884_),
    .A2(_10886_),
    .A3(_10889_),
    .S0(net518),
    .S1(net549),
    .X(_10892_));
 sky130_fd_sc_hd__mux2i_4 _25070_ (.A0(_10878_),
    .A1(_10892_),
    .S(net513),
    .Y(_10893_));
 sky130_fd_sc_hd__xnor2_1 _25071_ (.A(_10865_),
    .B(_10893_),
    .Y(_10894_));
 sky130_fd_sc_hd__xnor2_1 _25072_ (.A(_10833_),
    .B(_10894_),
    .Y(_11579_));
 sky130_fd_sc_hd__mux4_2 _25073_ (.A0(\w[1][4] ),
    .A1(\w[5][4] ),
    .A2(\w[3][4] ),
    .A3(\w[7][4] ),
    .S0(net521),
    .S1(net531),
    .X(_10895_));
 sky130_fd_sc_hd__mux4_2 _25074_ (.A0(\w[9][4] ),
    .A1(\w[13][4] ),
    .A2(\w[11][4] ),
    .A3(\w[15][4] ),
    .S0(net521),
    .S1(net531),
    .X(_10896_));
 sky130_fd_sc_hd__mux4_2 _25075_ (.A0(\w[17][4] ),
    .A1(\w[21][4] ),
    .A2(\w[19][4] ),
    .A3(\w[23][4] ),
    .S0(net521),
    .S1(net531),
    .X(_10897_));
 sky130_fd_sc_hd__mux4_2 _25076_ (.A0(\w[25][4] ),
    .A1(\w[29][4] ),
    .A2(\w[27][4] ),
    .A3(\w[31][4] ),
    .S0(net521),
    .S1(net531),
    .X(_10898_));
 sky130_fd_sc_hd__mux4_2 _25077_ (.A0(_10895_),
    .A1(_10896_),
    .A2(_10897_),
    .A3(_10898_),
    .S0(net516),
    .S1(net514),
    .X(_10899_));
 sky130_fd_sc_hd__mux4_2 _25078_ (.A0(\w[33][4] ),
    .A1(\w[37][4] ),
    .A2(\w[35][4] ),
    .A3(\w[39][4] ),
    .S0(net522),
    .S1(net531),
    .X(_10900_));
 sky130_fd_sc_hd__mux4_2 _25079_ (.A0(\w[41][4] ),
    .A1(\w[45][4] ),
    .A2(\w[43][4] ),
    .A3(\w[47][4] ),
    .S0(net522),
    .S1(net531),
    .X(_10901_));
 sky130_fd_sc_hd__mux4_2 _25080_ (.A0(\w[49][4] ),
    .A1(\w[53][4] ),
    .A2(\w[51][4] ),
    .A3(\w[55][4] ),
    .S0(net522),
    .S1(net531),
    .X(_10902_));
 sky130_fd_sc_hd__mux4_2 _25081_ (.A0(\w[57][4] ),
    .A1(\w[61][4] ),
    .A2(\w[59][4] ),
    .A3(\w[63][4] ),
    .S0(net522),
    .S1(net531),
    .X(_10903_));
 sky130_fd_sc_hd__mux4_2 _25082_ (.A0(_10900_),
    .A1(_10901_),
    .A2(_10902_),
    .A3(_10903_),
    .S0(net516),
    .S1(net514),
    .X(_10904_));
 sky130_fd_sc_hd__mux2i_4 _25083_ (.A0(_10899_),
    .A1(_10904_),
    .S(net512),
    .Y(_10905_));
 sky130_fd_sc_hd__mux4_2 _25084_ (.A0(\w[1][8] ),
    .A1(\w[5][8] ),
    .A2(\w[3][8] ),
    .A3(\w[7][8] ),
    .S0(net525),
    .S1(net529),
    .X(_10906_));
 sky130_fd_sc_hd__mux4_2 _25085_ (.A0(\w[9][8] ),
    .A1(\w[13][8] ),
    .A2(\w[11][8] ),
    .A3(\w[15][8] ),
    .S0(net525),
    .S1(net529),
    .X(_10907_));
 sky130_fd_sc_hd__mux4_2 _25086_ (.A0(\w[17][8] ),
    .A1(\w[21][8] ),
    .A2(\w[19][8] ),
    .A3(\w[23][8] ),
    .S0(net525),
    .S1(net529),
    .X(_10908_));
 sky130_fd_sc_hd__mux4_2 _25087_ (.A0(\w[25][8] ),
    .A1(\w[29][8] ),
    .A2(\w[27][8] ),
    .A3(\w[31][8] ),
    .S0(net525),
    .S1(net529),
    .X(_10909_));
 sky130_fd_sc_hd__mux4_2 _25088_ (.A0(_10906_),
    .A1(_10907_),
    .A2(_10908_),
    .A3(_10909_),
    .S0(net517),
    .S1(net514),
    .X(_10910_));
 sky130_fd_sc_hd__mux4_2 _25089_ (.A0(\w[33][8] ),
    .A1(\w[37][8] ),
    .A2(\w[35][8] ),
    .A3(\w[39][8] ),
    .S0(net526),
    .S1(net530),
    .X(_10911_));
 sky130_fd_sc_hd__mux4_2 _25090_ (.A0(\w[41][8] ),
    .A1(\w[45][8] ),
    .A2(\w[43][8] ),
    .A3(\w[47][8] ),
    .S0(net526),
    .S1(net530),
    .X(_10912_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_363 ();
 sky130_fd_sc_hd__mux4_2 _25092_ (.A0(\w[49][8] ),
    .A1(\w[53][8] ),
    .A2(\w[51][8] ),
    .A3(\w[55][8] ),
    .S0(net526),
    .S1(net530),
    .X(_10914_));
 sky130_fd_sc_hd__mux4_2 _25093_ (.A0(\w[57][8] ),
    .A1(\w[61][8] ),
    .A2(\w[59][8] ),
    .A3(\w[63][8] ),
    .S0(net526),
    .S1(net530),
    .X(_10915_));
 sky130_fd_sc_hd__mux4_2 _25094_ (.A0(_10911_),
    .A1(_10912_),
    .A2(_10914_),
    .A3(_10915_),
    .S0(net517),
    .S1(net514),
    .X(_10916_));
 sky130_fd_sc_hd__mux2i_4 _25095_ (.A0(_10910_),
    .A1(_10916_),
    .S(net512),
    .Y(_10917_));
 sky130_fd_sc_hd__mux4_2 _25096_ (.A0(\w[1][19] ),
    .A1(\w[5][19] ),
    .A2(\w[3][19] ),
    .A3(\w[7][19] ),
    .S0(net524),
    .S1(net529),
    .X(_10918_));
 sky130_fd_sc_hd__mux4_2 _25097_ (.A0(\w[9][19] ),
    .A1(\w[13][19] ),
    .A2(\w[11][19] ),
    .A3(\w[15][19] ),
    .S0(net524),
    .S1(net529),
    .X(_10919_));
 sky130_fd_sc_hd__mux4_2 _25098_ (.A0(\w[17][19] ),
    .A1(\w[21][19] ),
    .A2(\w[19][19] ),
    .A3(\w[23][19] ),
    .S0(net524),
    .S1(net529),
    .X(_10920_));
 sky130_fd_sc_hd__mux4_2 _25099_ (.A0(\w[25][19] ),
    .A1(\w[29][19] ),
    .A2(\w[27][19] ),
    .A3(\w[31][19] ),
    .S0(net524),
    .S1(net529),
    .X(_10921_));
 sky130_fd_sc_hd__mux4_2 _25100_ (.A0(_10918_),
    .A1(_10919_),
    .A2(_10920_),
    .A3(_10921_),
    .S0(net517),
    .S1(net515),
    .X(_10922_));
 sky130_fd_sc_hd__mux4_2 _25101_ (.A0(\w[33][19] ),
    .A1(\w[37][19] ),
    .A2(\w[35][19] ),
    .A3(\w[39][19] ),
    .S0(net527),
    .S1(net550),
    .X(_10923_));
 sky130_fd_sc_hd__mux4_2 _25102_ (.A0(\w[41][19] ),
    .A1(\w[45][19] ),
    .A2(\w[43][19] ),
    .A3(\w[47][19] ),
    .S0(net527),
    .S1(net550),
    .X(_10924_));
 sky130_fd_sc_hd__mux4_2 _25103_ (.A0(\w[49][19] ),
    .A1(\w[53][19] ),
    .A2(\w[51][19] ),
    .A3(\w[55][19] ),
    .S0(net527),
    .S1(net550),
    .X(_10925_));
 sky130_fd_sc_hd__mux4_2 _25104_ (.A0(\w[57][19] ),
    .A1(\w[61][19] ),
    .A2(\w[59][19] ),
    .A3(\w[63][19] ),
    .S0(net527),
    .S1(net550),
    .X(_10926_));
 sky130_fd_sc_hd__mux4_2 _25105_ (.A0(_10923_),
    .A1(_10924_),
    .A2(_10925_),
    .A3(_10926_),
    .S0(\count15_1[3] ),
    .S1(net515),
    .X(_10927_));
 sky130_fd_sc_hd__mux2i_4 _25106_ (.A0(_10922_),
    .A1(_10927_),
    .S(\count15_1[5] ),
    .Y(_10928_));
 sky130_fd_sc_hd__xnor2_1 _25107_ (.A(_10917_),
    .B(_10928_),
    .Y(_10929_));
 sky130_fd_sc_hd__xnor2_1 _25108_ (.A(_10905_),
    .B(_10929_),
    .Y(_11584_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_353 ();
 sky130_fd_sc_hd__mux4_2 _25119_ (.A0(\w[0][11] ),
    .A1(\w[4][11] ),
    .A2(\w[2][11] ),
    .A3(\w[6][11] ),
    .S0(net442),
    .S1(net450),
    .X(_10940_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_351 ();
 sky130_fd_sc_hd__mux4_2 _25122_ (.A0(\w[8][11] ),
    .A1(\w[12][11] ),
    .A2(\w[10][11] ),
    .A3(\w[14][11] ),
    .S0(net442),
    .S1(net450),
    .X(_10943_));
 sky130_fd_sc_hd__mux4_2 _25123_ (.A0(\w[16][11] ),
    .A1(\w[20][11] ),
    .A2(\w[18][11] ),
    .A3(\w[22][11] ),
    .S0(net440),
    .S1(net448),
    .X(_10944_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_349 ();
 sky130_fd_sc_hd__mux4_2 _25126_ (.A0(\w[24][11] ),
    .A1(\w[28][11] ),
    .A2(\w[26][11] ),
    .A3(\w[30][11] ),
    .S0(net440),
    .S1(net448),
    .X(_10947_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_344 ();
 sky130_fd_sc_hd__mux4_2 _25132_ (.A0(_10940_),
    .A1(_10943_),
    .A2(_10944_),
    .A3(_10947_),
    .S0(net438),
    .S1(net434),
    .X(_10953_));
 sky130_fd_sc_hd__mux4_2 _25133_ (.A0(\w[32][11] ),
    .A1(\w[36][11] ),
    .A2(\w[34][11] ),
    .A3(\w[38][11] ),
    .S0(net443),
    .S1(net451),
    .X(_10954_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_342 ();
 sky130_fd_sc_hd__mux4_2 _25136_ (.A0(\w[40][11] ),
    .A1(\w[44][11] ),
    .A2(\w[42][11] ),
    .A3(\w[46][11] ),
    .S0(net443),
    .S1(net451),
    .X(_10957_));
 sky130_fd_sc_hd__mux4_2 _25137_ (.A0(\w[48][11] ),
    .A1(\w[52][11] ),
    .A2(\w[50][11] ),
    .A3(\w[54][11] ),
    .S0(net443),
    .S1(net451),
    .X(_10958_));
 sky130_fd_sc_hd__mux4_2 _25138_ (.A0(\w[56][11] ),
    .A1(\w[60][11] ),
    .A2(\w[58][11] ),
    .A3(\w[62][11] ),
    .S0(net443),
    .S1(net451),
    .X(_10959_));
 sky130_fd_sc_hd__mux4_2 _25139_ (.A0(_10954_),
    .A1(_10957_),
    .A2(_10958_),
    .A3(_10959_),
    .S0(net436),
    .S1(net434),
    .X(_10960_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_340 ();
 sky130_fd_sc_hd__mux2i_4 _25142_ (.A0(_10953_),
    .A1(_10960_),
    .S(net432),
    .Y(_10963_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_337 ();
 sky130_fd_sc_hd__mux4_2 _25146_ (.A0(\w[0][20] ),
    .A1(\w[4][20] ),
    .A2(\w[2][20] ),
    .A3(\w[6][20] ),
    .S0(net441),
    .S1(net449),
    .X(_10967_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_335 ();
 sky130_fd_sc_hd__mux4_2 _25149_ (.A0(\w[8][20] ),
    .A1(\w[12][20] ),
    .A2(\w[10][20] ),
    .A3(\w[14][20] ),
    .S0(net441),
    .S1(net449),
    .X(_10970_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_333 ();
 sky130_fd_sc_hd__mux4_2 _25152_ (.A0(\w[16][20] ),
    .A1(\w[20][20] ),
    .A2(\w[18][20] ),
    .A3(\w[22][20] ),
    .S0(net441),
    .S1(net449),
    .X(_10973_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_331 ();
 sky130_fd_sc_hd__mux4_2 _25155_ (.A0(\w[24][20] ),
    .A1(\w[28][20] ),
    .A2(\w[26][20] ),
    .A3(\w[30][20] ),
    .S0(net441),
    .S1(net449),
    .X(_10976_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_329 ();
 sky130_fd_sc_hd__mux4_2 _25158_ (.A0(_10967_),
    .A1(_10970_),
    .A2(_10973_),
    .A3(_10976_),
    .S0(net436),
    .S1(net434),
    .X(_10979_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_327 ();
 sky130_fd_sc_hd__mux4_2 _25161_ (.A0(\w[32][20] ),
    .A1(\w[36][20] ),
    .A2(\w[34][20] ),
    .A3(\w[38][20] ),
    .S0(net443),
    .S1(net451),
    .X(_10982_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_326 ();
 sky130_fd_sc_hd__mux4_2 _25163_ (.A0(\w[40][20] ),
    .A1(\w[44][20] ),
    .A2(\w[42][20] ),
    .A3(\w[46][20] ),
    .S0(net443),
    .S1(net451),
    .X(_10984_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_324 ();
 sky130_fd_sc_hd__mux4_2 _25166_ (.A0(\w[48][20] ),
    .A1(\w[52][20] ),
    .A2(\w[50][20] ),
    .A3(\w[54][20] ),
    .S0(net443),
    .S1(net451),
    .X(_10987_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_322 ();
 sky130_fd_sc_hd__mux4_2 _25169_ (.A0(\w[56][20] ),
    .A1(\w[60][20] ),
    .A2(\w[58][20] ),
    .A3(\w[62][20] ),
    .S0(net443),
    .S1(net451),
    .X(_10990_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_320 ();
 sky130_fd_sc_hd__mux4_2 _25172_ (.A0(_10982_),
    .A1(_10984_),
    .A2(_10987_),
    .A3(_10990_),
    .S0(net436),
    .S1(net434),
    .X(_10993_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_319 ();
 sky130_fd_sc_hd__mux2i_4 _25174_ (.A0(_10979_),
    .A1(_10993_),
    .S(net432),
    .Y(_10995_));
 sky130_fd_sc_hd__mux4_2 _25175_ (.A0(\w[0][18] ),
    .A1(\w[4][18] ),
    .A2(\w[2][18] ),
    .A3(\w[6][18] ),
    .S0(net443),
    .S1(net451),
    .X(_10996_));
 sky130_fd_sc_hd__mux4_2 _25176_ (.A0(\w[8][18] ),
    .A1(\w[12][18] ),
    .A2(\w[10][18] ),
    .A3(\w[14][18] ),
    .S0(net443),
    .S1(net451),
    .X(_10997_));
 sky130_fd_sc_hd__mux4_2 _25177_ (.A0(\w[16][18] ),
    .A1(\w[20][18] ),
    .A2(\w[18][18] ),
    .A3(\w[22][18] ),
    .S0(net443),
    .S1(net451),
    .X(_10998_));
 sky130_fd_sc_hd__mux4_2 _25178_ (.A0(\w[24][18] ),
    .A1(\w[28][18] ),
    .A2(\w[26][18] ),
    .A3(\w[30][18] ),
    .S0(net443),
    .S1(net451),
    .X(_10999_));
 sky130_fd_sc_hd__mux4_2 _25179_ (.A0(_10996_),
    .A1(_10997_),
    .A2(_10998_),
    .A3(_10999_),
    .S0(net436),
    .S1(net434),
    .X(_11000_));
 sky130_fd_sc_hd__mux4_2 _25180_ (.A0(\w[32][18] ),
    .A1(\w[36][18] ),
    .A2(\w[34][18] ),
    .A3(\w[38][18] ),
    .S0(net443),
    .S1(net451),
    .X(_11001_));
 sky130_fd_sc_hd__mux4_2 _25181_ (.A0(\w[40][18] ),
    .A1(\w[44][18] ),
    .A2(\w[42][18] ),
    .A3(\w[46][18] ),
    .S0(net443),
    .S1(net451),
    .X(_11002_));
 sky130_fd_sc_hd__mux4_2 _25182_ (.A0(\w[48][18] ),
    .A1(\w[52][18] ),
    .A2(\w[50][18] ),
    .A3(\w[54][18] ),
    .S0(net443),
    .S1(net451),
    .X(_11003_));
 sky130_fd_sc_hd__mux4_2 _25183_ (.A0(\w[56][18] ),
    .A1(\w[60][18] ),
    .A2(\w[58][18] ),
    .A3(\w[62][18] ),
    .S0(net443),
    .S1(net451),
    .X(_11004_));
 sky130_fd_sc_hd__mux4_2 _25184_ (.A0(_11001_),
    .A1(_11002_),
    .A2(_11003_),
    .A3(_11004_),
    .S0(net436),
    .S1(net434),
    .X(_11005_));
 sky130_fd_sc_hd__mux2i_4 _25185_ (.A0(_11000_),
    .A1(_11005_),
    .S(net432),
    .Y(_11006_));
 sky130_fd_sc_hd__xnor2_1 _25186_ (.A(_10995_),
    .B(_11006_),
    .Y(_11007_));
 sky130_fd_sc_hd__xnor2_1 _25187_ (.A(_10963_),
    .B(_11007_),
    .Y(_11589_));
 sky130_fd_sc_hd__mux4_2 _25188_ (.A0(\w[1][20] ),
    .A1(\w[5][20] ),
    .A2(\w[3][20] ),
    .A3(\w[7][20] ),
    .S0(net524),
    .S1(net530),
    .X(_11008_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_318 ();
 sky130_fd_sc_hd__mux4_2 _25190_ (.A0(\w[9][20] ),
    .A1(\w[13][20] ),
    .A2(\w[11][20] ),
    .A3(\w[15][20] ),
    .S0(net524),
    .S1(net530),
    .X(_11010_));
 sky130_fd_sc_hd__mux4_2 _25191_ (.A0(\w[17][20] ),
    .A1(\w[21][20] ),
    .A2(\w[19][20] ),
    .A3(\w[23][20] ),
    .S0(net524),
    .S1(net530),
    .X(_11011_));
 sky130_fd_sc_hd__mux4_2 _25192_ (.A0(\w[25][20] ),
    .A1(\w[29][20] ),
    .A2(\w[27][20] ),
    .A3(\w[31][20] ),
    .S0(net524),
    .S1(net530),
    .X(_11012_));
 sky130_fd_sc_hd__mux4_2 _25193_ (.A0(_11008_),
    .A1(_11010_),
    .A2(_11011_),
    .A3(_11012_),
    .S0(net517),
    .S1(net515),
    .X(_11013_));
 sky130_fd_sc_hd__mux4_2 _25194_ (.A0(\w[33][20] ),
    .A1(\w[37][20] ),
    .A2(\w[35][20] ),
    .A3(\w[39][20] ),
    .S0(net527),
    .S1(net550),
    .X(_11014_));
 sky130_fd_sc_hd__mux4_2 _25195_ (.A0(\w[41][20] ),
    .A1(\w[45][20] ),
    .A2(\w[43][20] ),
    .A3(\w[47][20] ),
    .S0(net527),
    .S1(net550),
    .X(_11015_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_317 ();
 sky130_fd_sc_hd__mux4_2 _25197_ (.A0(\w[49][20] ),
    .A1(\w[53][20] ),
    .A2(\w[51][20] ),
    .A3(\w[55][20] ),
    .S0(net527),
    .S1(net550),
    .X(_11017_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_315 ();
 sky130_fd_sc_hd__mux4_2 _25200_ (.A0(\w[57][20] ),
    .A1(\w[61][20] ),
    .A2(\w[59][20] ),
    .A3(\w[63][20] ),
    .S0(net527),
    .S1(net550),
    .X(_11020_));
 sky130_fd_sc_hd__mux4_2 _25201_ (.A0(_11014_),
    .A1(_11015_),
    .A2(_11017_),
    .A3(_11020_),
    .S0(\count15_1[3] ),
    .S1(net515),
    .X(_11021_));
 sky130_fd_sc_hd__mux2i_4 _25202_ (.A0(_11013_),
    .A1(_11021_),
    .S(\count15_1[5] ),
    .Y(_11022_));
 sky130_fd_sc_hd__mux4_2 _25203_ (.A0(\w[1][5] ),
    .A1(\w[5][5] ),
    .A2(\w[3][5] ),
    .A3(\w[7][5] ),
    .S0(net519),
    .S1(net528),
    .X(_11023_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_314 ();
 sky130_fd_sc_hd__mux4_2 _25205_ (.A0(\w[9][5] ),
    .A1(\w[13][5] ),
    .A2(\w[11][5] ),
    .A3(\w[15][5] ),
    .S0(net519),
    .S1(net528),
    .X(_11025_));
 sky130_fd_sc_hd__mux4_2 _25206_ (.A0(\w[17][5] ),
    .A1(\w[21][5] ),
    .A2(\w[19][5] ),
    .A3(\w[23][5] ),
    .S0(net519),
    .S1(net528),
    .X(_11026_));
 sky130_fd_sc_hd__mux4_2 _25207_ (.A0(\w[25][5] ),
    .A1(\w[29][5] ),
    .A2(\w[27][5] ),
    .A3(\w[31][5] ),
    .S0(net519),
    .S1(net528),
    .X(_11027_));
 sky130_fd_sc_hd__mux4_2 _25208_ (.A0(_11023_),
    .A1(_11025_),
    .A2(_11026_),
    .A3(_11027_),
    .S0(net516),
    .S1(net514),
    .X(_11028_));
 sky130_fd_sc_hd__mux4_2 _25209_ (.A0(\w[33][5] ),
    .A1(\w[37][5] ),
    .A2(\w[35][5] ),
    .A3(\w[39][5] ),
    .S0(net519),
    .S1(net528),
    .X(_11029_));
 sky130_fd_sc_hd__mux4_2 _25210_ (.A0(\w[41][5] ),
    .A1(\w[45][5] ),
    .A2(\w[43][5] ),
    .A3(\w[47][5] ),
    .S0(net519),
    .S1(net528),
    .X(_11030_));
 sky130_fd_sc_hd__mux4_2 _25211_ (.A0(\w[49][5] ),
    .A1(\w[53][5] ),
    .A2(\w[51][5] ),
    .A3(\w[55][5] ),
    .S0(net519),
    .S1(net528),
    .X(_11031_));
 sky130_fd_sc_hd__mux4_2 _25212_ (.A0(\w[57][5] ),
    .A1(\w[61][5] ),
    .A2(\w[59][5] ),
    .A3(\w[63][5] ),
    .S0(net519),
    .S1(net528),
    .X(_11032_));
 sky130_fd_sc_hd__mux4_2 _25213_ (.A0(_11029_),
    .A1(_11030_),
    .A2(_11031_),
    .A3(_11032_),
    .S0(net518),
    .S1(net549),
    .X(_11033_));
 sky130_fd_sc_hd__mux2i_4 _25214_ (.A0(_11028_),
    .A1(_11033_),
    .S(net513),
    .Y(_11034_));
 sky130_fd_sc_hd__mux4_2 _25215_ (.A0(\w[1][9] ),
    .A1(\w[5][9] ),
    .A2(\w[3][9] ),
    .A3(\w[7][9] ),
    .S0(net523),
    .S1(net532),
    .X(_11035_));
 sky130_fd_sc_hd__mux4_2 _25216_ (.A0(\w[9][9] ),
    .A1(\w[13][9] ),
    .A2(\w[11][9] ),
    .A3(\w[15][9] ),
    .S0(net523),
    .S1(net532),
    .X(_11036_));
 sky130_fd_sc_hd__mux4_2 _25217_ (.A0(\w[17][9] ),
    .A1(\w[21][9] ),
    .A2(\w[19][9] ),
    .A3(\w[23][9] ),
    .S0(net523),
    .S1(net532),
    .X(_11037_));
 sky130_fd_sc_hd__mux4_2 _25218_ (.A0(\w[25][9] ),
    .A1(\w[29][9] ),
    .A2(\w[27][9] ),
    .A3(\w[31][9] ),
    .S0(net523),
    .S1(net532),
    .X(_11038_));
 sky130_fd_sc_hd__mux4_2 _25219_ (.A0(_11035_),
    .A1(_11036_),
    .A2(_11037_),
    .A3(_11038_),
    .S0(net518),
    .S1(net549),
    .X(_11039_));
 sky130_fd_sc_hd__mux4_2 _25220_ (.A0(\w[33][9] ),
    .A1(\w[37][9] ),
    .A2(\w[35][9] ),
    .A3(\w[39][9] ),
    .S0(net522),
    .S1(\count15_1[1] ),
    .X(_11040_));
 sky130_fd_sc_hd__mux4_2 _25221_ (.A0(\w[41][9] ),
    .A1(\w[45][9] ),
    .A2(\w[43][9] ),
    .A3(\w[47][9] ),
    .S0(net522),
    .S1(\count15_1[1] ),
    .X(_11041_));
 sky130_fd_sc_hd__mux4_2 _25222_ (.A0(\w[49][9] ),
    .A1(\w[53][9] ),
    .A2(\w[51][9] ),
    .A3(\w[55][9] ),
    .S0(net522),
    .S1(\count15_1[1] ),
    .X(_11042_));
 sky130_fd_sc_hd__mux4_2 _25223_ (.A0(\w[57][9] ),
    .A1(\w[61][9] ),
    .A2(\w[59][9] ),
    .A3(\w[63][9] ),
    .S0(net522),
    .S1(\count15_1[1] ),
    .X(_11043_));
 sky130_fd_sc_hd__mux4_2 _25224_ (.A0(_11040_),
    .A1(_11041_),
    .A2(_11042_),
    .A3(_11043_),
    .S0(net516),
    .S1(net514),
    .X(_11044_));
 sky130_fd_sc_hd__mux2i_4 _25225_ (.A0(_11039_),
    .A1(_11044_),
    .S(net513),
    .Y(_11045_));
 sky130_fd_sc_hd__xnor2_1 _25226_ (.A(_11034_),
    .B(_11045_),
    .Y(_11046_));
 sky130_fd_sc_hd__xnor2_1 _25227_ (.A(_11022_),
    .B(_11046_),
    .Y(_11592_));
 sky130_fd_sc_hd__mux4_2 _25228_ (.A0(\w[0][12] ),
    .A1(\w[4][12] ),
    .A2(\w[2][12] ),
    .A3(\w[6][12] ),
    .S0(net445),
    .S1(net452),
    .X(_11047_));
 sky130_fd_sc_hd__mux4_2 _25229_ (.A0(\w[8][12] ),
    .A1(\w[12][12] ),
    .A2(\w[10][12] ),
    .A3(\w[14][12] ),
    .S0(net445),
    .S1(net452),
    .X(_11048_));
 sky130_fd_sc_hd__mux4_2 _25230_ (.A0(\w[16][12] ),
    .A1(\w[20][12] ),
    .A2(\w[18][12] ),
    .A3(\w[22][12] ),
    .S0(net445),
    .S1(net452),
    .X(_11049_));
 sky130_fd_sc_hd__mux4_2 _25231_ (.A0(\w[24][12] ),
    .A1(\w[28][12] ),
    .A2(\w[26][12] ),
    .A3(\w[30][12] ),
    .S0(net445),
    .S1(net452),
    .X(_11050_));
 sky130_fd_sc_hd__mux4_2 _25232_ (.A0(_11047_),
    .A1(_11048_),
    .A2(_11049_),
    .A3(_11050_),
    .S0(net437),
    .S1(net435),
    .X(_11051_));
 sky130_fd_sc_hd__mux4_2 _25233_ (.A0(\w[32][12] ),
    .A1(\w[36][12] ),
    .A2(\w[34][12] ),
    .A3(\w[38][12] ),
    .S0(net445),
    .S1(net452),
    .X(_11052_));
 sky130_fd_sc_hd__mux4_2 _25234_ (.A0(\w[40][12] ),
    .A1(\w[44][12] ),
    .A2(\w[42][12] ),
    .A3(\w[46][12] ),
    .S0(net445),
    .S1(net452),
    .X(_11053_));
 sky130_fd_sc_hd__mux4_2 _25235_ (.A0(\w[48][12] ),
    .A1(\w[52][12] ),
    .A2(\w[50][12] ),
    .A3(\w[54][12] ),
    .S0(net445),
    .S1(net452),
    .X(_11054_));
 sky130_fd_sc_hd__mux4_2 _25236_ (.A0(\w[56][12] ),
    .A1(\w[60][12] ),
    .A2(\w[58][12] ),
    .A3(\w[62][12] ),
    .S0(net445),
    .S1(net452),
    .X(_11055_));
 sky130_fd_sc_hd__mux4_2 _25237_ (.A0(_11052_),
    .A1(_11053_),
    .A2(_11054_),
    .A3(_11055_),
    .S0(net437),
    .S1(net435),
    .X(_11056_));
 sky130_fd_sc_hd__mux2i_4 _25238_ (.A0(_11051_),
    .A1(_11056_),
    .S(net433),
    .Y(_11057_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_313 ();
 sky130_fd_sc_hd__mux4_2 _25240_ (.A0(\w[0][21] ),
    .A1(\w[4][21] ),
    .A2(\w[2][21] ),
    .A3(\w[6][21] ),
    .S0(net440),
    .S1(net448),
    .X(_11059_));
 sky130_fd_sc_hd__mux4_2 _25241_ (.A0(\w[8][21] ),
    .A1(\w[12][21] ),
    .A2(\w[10][21] ),
    .A3(\w[14][21] ),
    .S0(net440),
    .S1(net448),
    .X(_11060_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_312 ();
 sky130_fd_sc_hd__mux4_2 _25243_ (.A0(\w[16][21] ),
    .A1(\w[20][21] ),
    .A2(\w[18][21] ),
    .A3(\w[22][21] ),
    .S0(net440),
    .S1(net448),
    .X(_11062_));
 sky130_fd_sc_hd__mux4_2 _25244_ (.A0(\w[24][21] ),
    .A1(\w[28][21] ),
    .A2(\w[26][21] ),
    .A3(\w[30][21] ),
    .S0(net440),
    .S1(net448),
    .X(_11063_));
 sky130_fd_sc_hd__mux4_2 _25245_ (.A0(_11059_),
    .A1(_11060_),
    .A2(_11062_),
    .A3(_11063_),
    .S0(net438),
    .S1(net434),
    .X(_11064_));
 sky130_fd_sc_hd__mux4_2 _25246_ (.A0(\w[32][21] ),
    .A1(\w[36][21] ),
    .A2(\w[34][21] ),
    .A3(\w[38][21] ),
    .S0(net443),
    .S1(net451),
    .X(_11065_));
 sky130_fd_sc_hd__mux4_2 _25247_ (.A0(\w[40][21] ),
    .A1(\w[44][21] ),
    .A2(\w[42][21] ),
    .A3(\w[46][21] ),
    .S0(net443),
    .S1(net451),
    .X(_11066_));
 sky130_fd_sc_hd__mux4_2 _25248_ (.A0(\w[48][21] ),
    .A1(\w[52][21] ),
    .A2(\w[50][21] ),
    .A3(\w[54][21] ),
    .S0(net443),
    .S1(net451),
    .X(_11067_));
 sky130_fd_sc_hd__mux4_2 _25249_ (.A0(\w[56][21] ),
    .A1(\w[60][21] ),
    .A2(\w[58][21] ),
    .A3(\w[62][21] ),
    .S0(net443),
    .S1(net451),
    .X(_11068_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_311 ();
 sky130_fd_sc_hd__mux4_2 _25251_ (.A0(_11065_),
    .A1(_11066_),
    .A2(_11067_),
    .A3(_11068_),
    .S0(net436),
    .S1(net434),
    .X(_11070_));
 sky130_fd_sc_hd__mux2i_4 _25252_ (.A0(_11064_),
    .A1(_11070_),
    .S(net432),
    .Y(_11071_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_310 ();
 sky130_fd_sc_hd__mux4_2 _25254_ (.A0(\w[0][19] ),
    .A1(\w[4][19] ),
    .A2(\w[2][19] ),
    .A3(\w[6][19] ),
    .S0(net440),
    .S1(net448),
    .X(_11073_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_309 ();
 sky130_fd_sc_hd__mux4_2 _25256_ (.A0(\w[8][19] ),
    .A1(\w[12][19] ),
    .A2(\w[10][19] ),
    .A3(\w[14][19] ),
    .S0(net440),
    .S1(net448),
    .X(_11075_));
 sky130_fd_sc_hd__mux4_2 _25257_ (.A0(\w[16][19] ),
    .A1(\w[20][19] ),
    .A2(\w[18][19] ),
    .A3(\w[22][19] ),
    .S0(net440),
    .S1(net448),
    .X(_11076_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_307 ();
 sky130_fd_sc_hd__mux4_2 _25260_ (.A0(\w[24][19] ),
    .A1(\w[28][19] ),
    .A2(\w[26][19] ),
    .A3(\w[30][19] ),
    .S0(net440),
    .S1(net448),
    .X(_11079_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_305 ();
 sky130_fd_sc_hd__mux4_2 _25263_ (.A0(_11073_),
    .A1(_11075_),
    .A2(_11076_),
    .A3(_11079_),
    .S0(net438),
    .S1(net434),
    .X(_11082_));
 sky130_fd_sc_hd__mux4_2 _25264_ (.A0(\w[32][19] ),
    .A1(\w[36][19] ),
    .A2(\w[34][19] ),
    .A3(\w[38][19] ),
    .S0(net441),
    .S1(net449),
    .X(_11083_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_303 ();
 sky130_fd_sc_hd__mux4_2 _25267_ (.A0(\w[40][19] ),
    .A1(\w[44][19] ),
    .A2(\w[42][19] ),
    .A3(\w[46][19] ),
    .S0(net441),
    .S1(net449),
    .X(_11086_));
 sky130_fd_sc_hd__mux4_2 _25268_ (.A0(\w[48][19] ),
    .A1(\w[52][19] ),
    .A2(\w[50][19] ),
    .A3(\w[54][19] ),
    .S0(net441),
    .S1(net449),
    .X(_11087_));
 sky130_fd_sc_hd__mux4_2 _25269_ (.A0(\w[56][19] ),
    .A1(\w[60][19] ),
    .A2(\w[58][19] ),
    .A3(\w[62][19] ),
    .S0(net441),
    .S1(net449),
    .X(_11088_));
 sky130_fd_sc_hd__mux4_2 _25270_ (.A0(_11083_),
    .A1(_11086_),
    .A2(_11087_),
    .A3(_11088_),
    .S0(net436),
    .S1(net434),
    .X(_11089_));
 sky130_fd_sc_hd__mux2i_4 _25271_ (.A0(_11082_),
    .A1(_11089_),
    .S(net432),
    .Y(_11090_));
 sky130_fd_sc_hd__xnor2_1 _25272_ (.A(_11071_),
    .B(_11090_),
    .Y(_11091_));
 sky130_fd_sc_hd__xnor2_1 _25273_ (.A(_11057_),
    .B(_11091_),
    .Y(_11597_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_301 ();
 sky130_fd_sc_hd__mux4_2 _25276_ (.A0(\w[1][6] ),
    .A1(\w[5][6] ),
    .A2(\w[3][6] ),
    .A3(\w[7][6] ),
    .S0(net526),
    .S1(net529),
    .X(_11094_));
 sky130_fd_sc_hd__mux4_2 _25277_ (.A0(\w[9][6] ),
    .A1(\w[13][6] ),
    .A2(\w[11][6] ),
    .A3(\w[15][6] ),
    .S0(net526),
    .S1(net529),
    .X(_11095_));
 sky130_fd_sc_hd__mux4_2 _25278_ (.A0(\w[17][6] ),
    .A1(\w[21][6] ),
    .A2(\w[19][6] ),
    .A3(\w[23][6] ),
    .S0(net526),
    .S1(net529),
    .X(_11096_));
 sky130_fd_sc_hd__mux4_2 _25279_ (.A0(\w[25][6] ),
    .A1(\w[29][6] ),
    .A2(\w[27][6] ),
    .A3(\w[31][6] ),
    .S0(net526),
    .S1(net529),
    .X(_11097_));
 sky130_fd_sc_hd__mux4_2 _25280_ (.A0(_11094_),
    .A1(_11095_),
    .A2(_11096_),
    .A3(_11097_),
    .S0(net517),
    .S1(net514),
    .X(_11098_));
 sky130_fd_sc_hd__mux4_2 _25281_ (.A0(\w[33][6] ),
    .A1(\w[37][6] ),
    .A2(\w[35][6] ),
    .A3(\w[39][6] ),
    .S0(net526),
    .S1(net530),
    .X(_11099_));
 sky130_fd_sc_hd__mux4_2 _25282_ (.A0(\w[41][6] ),
    .A1(\w[45][6] ),
    .A2(\w[43][6] ),
    .A3(\w[47][6] ),
    .S0(net526),
    .S1(net530),
    .X(_11100_));
 sky130_fd_sc_hd__mux4_2 _25283_ (.A0(\w[49][6] ),
    .A1(\w[53][6] ),
    .A2(\w[51][6] ),
    .A3(\w[55][6] ),
    .S0(net526),
    .S1(net530),
    .X(_11101_));
 sky130_fd_sc_hd__mux4_2 _25284_ (.A0(\w[57][6] ),
    .A1(\w[61][6] ),
    .A2(\w[59][6] ),
    .A3(\w[63][6] ),
    .S0(net526),
    .S1(net530),
    .X(_11102_));
 sky130_fd_sc_hd__mux4_2 _25285_ (.A0(_11099_),
    .A1(_11100_),
    .A2(_11101_),
    .A3(_11102_),
    .S0(net517),
    .S1(net514),
    .X(_11103_));
 sky130_fd_sc_hd__mux2i_4 _25286_ (.A0(_11098_),
    .A1(_11103_),
    .S(net512),
    .Y(_11104_));
 sky130_fd_sc_hd__mux4_2 _25287_ (.A0(\w[1][21] ),
    .A1(\w[5][21] ),
    .A2(\w[3][21] ),
    .A3(\w[7][21] ),
    .S0(net524),
    .S1(net529),
    .X(_11105_));
 sky130_fd_sc_hd__mux4_2 _25288_ (.A0(\w[9][21] ),
    .A1(\w[13][21] ),
    .A2(\w[11][21] ),
    .A3(\w[15][21] ),
    .S0(net524),
    .S1(net529),
    .X(_11106_));
 sky130_fd_sc_hd__mux4_2 _25289_ (.A0(\w[17][21] ),
    .A1(\w[21][21] ),
    .A2(\w[19][21] ),
    .A3(\w[23][21] ),
    .S0(net524),
    .S1(net529),
    .X(_11107_));
 sky130_fd_sc_hd__mux4_2 _25290_ (.A0(\w[25][21] ),
    .A1(\w[29][21] ),
    .A2(\w[27][21] ),
    .A3(\w[31][21] ),
    .S0(net524),
    .S1(net529),
    .X(_11108_));
 sky130_fd_sc_hd__mux4_2 _25291_ (.A0(_11105_),
    .A1(_11106_),
    .A2(_11107_),
    .A3(_11108_),
    .S0(net517),
    .S1(net515),
    .X(_11109_));
 sky130_fd_sc_hd__mux4_2 _25292_ (.A0(\w[33][21] ),
    .A1(\w[37][21] ),
    .A2(\w[35][21] ),
    .A3(\w[39][21] ),
    .S0(net525),
    .S1(net530),
    .X(_11110_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_300 ();
 sky130_fd_sc_hd__mux4_2 _25294_ (.A0(\w[41][21] ),
    .A1(\w[45][21] ),
    .A2(\w[43][21] ),
    .A3(\w[47][21] ),
    .S0(net525),
    .S1(net530),
    .X(_11112_));
 sky130_fd_sc_hd__mux4_2 _25295_ (.A0(\w[49][21] ),
    .A1(\w[53][21] ),
    .A2(\w[51][21] ),
    .A3(\w[55][21] ),
    .S0(net525),
    .S1(net530),
    .X(_11113_));
 sky130_fd_sc_hd__mux4_2 _25296_ (.A0(\w[57][21] ),
    .A1(\w[61][21] ),
    .A2(\w[59][21] ),
    .A3(\w[63][21] ),
    .S0(net525),
    .S1(net530),
    .X(_11114_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_299 ();
 sky130_fd_sc_hd__mux4_2 _25298_ (.A0(_11110_),
    .A1(_11112_),
    .A2(_11113_),
    .A3(_11114_),
    .S0(net517),
    .S1(net515),
    .X(_11116_));
 sky130_fd_sc_hd__mux2i_4 _25299_ (.A0(_11109_),
    .A1(_11116_),
    .S(\count15_1[5] ),
    .Y(_11117_));
 sky130_fd_sc_hd__mux4_2 _25300_ (.A0(\w[1][10] ),
    .A1(\w[5][10] ),
    .A2(\w[3][10] ),
    .A3(\w[7][10] ),
    .S0(net524),
    .S1(net530),
    .X(_11118_));
 sky130_fd_sc_hd__mux4_2 _25301_ (.A0(\w[9][10] ),
    .A1(\w[13][10] ),
    .A2(\w[11][10] ),
    .A3(\w[15][10] ),
    .S0(net524),
    .S1(net530),
    .X(_11119_));
 sky130_fd_sc_hd__mux4_2 _25302_ (.A0(\w[17][10] ),
    .A1(\w[21][10] ),
    .A2(\w[19][10] ),
    .A3(\w[23][10] ),
    .S0(net524),
    .S1(net530),
    .X(_11120_));
 sky130_fd_sc_hd__mux4_2 _25303_ (.A0(\w[25][10] ),
    .A1(\w[29][10] ),
    .A2(\w[27][10] ),
    .A3(\w[31][10] ),
    .S0(net524),
    .S1(net530),
    .X(_11121_));
 sky130_fd_sc_hd__mux4_2 _25304_ (.A0(_11118_),
    .A1(_11119_),
    .A2(_11120_),
    .A3(_11121_),
    .S0(net517),
    .S1(net515),
    .X(_11122_));
 sky130_fd_sc_hd__mux4_2 _25305_ (.A0(\w[33][10] ),
    .A1(\w[37][10] ),
    .A2(\w[35][10] ),
    .A3(\w[39][10] ),
    .S0(net525),
    .S1(net530),
    .X(_11123_));
 sky130_fd_sc_hd__mux4_2 _25306_ (.A0(\w[41][10] ),
    .A1(\w[45][10] ),
    .A2(\w[43][10] ),
    .A3(\w[47][10] ),
    .S0(net525),
    .S1(net530),
    .X(_11124_));
 sky130_fd_sc_hd__mux4_2 _25307_ (.A0(\w[49][10] ),
    .A1(\w[53][10] ),
    .A2(\w[51][10] ),
    .A3(\w[55][10] ),
    .S0(net526),
    .S1(net530),
    .X(_11125_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_298 ();
 sky130_fd_sc_hd__mux4_2 _25309_ (.A0(\w[57][10] ),
    .A1(\w[61][10] ),
    .A2(\w[59][10] ),
    .A3(\w[63][10] ),
    .S0(net526),
    .S1(net530),
    .X(_11127_));
 sky130_fd_sc_hd__mux4_2 _25310_ (.A0(_11123_),
    .A1(_11124_),
    .A2(_11125_),
    .A3(_11127_),
    .S0(net517),
    .S1(net515),
    .X(_11128_));
 sky130_fd_sc_hd__mux2i_4 _25311_ (.A0(_11122_),
    .A1(_11128_),
    .S(\count15_1[5] ),
    .Y(_11129_));
 sky130_fd_sc_hd__xnor2_1 _25312_ (.A(_11117_),
    .B(_11129_),
    .Y(_11130_));
 sky130_fd_sc_hd__xnor2_1 _25313_ (.A(_11104_),
    .B(_11130_),
    .Y(_11603_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_297 ();
 sky130_fd_sc_hd__mux4_2 _25315_ (.A0(\w[0][13] ),
    .A1(\w[4][13] ),
    .A2(\w[2][13] ),
    .A3(\w[6][13] ),
    .S0(net442),
    .S1(net450),
    .X(_11132_));
 sky130_fd_sc_hd__mux4_2 _25316_ (.A0(\w[8][13] ),
    .A1(\w[12][13] ),
    .A2(\w[10][13] ),
    .A3(\w[14][13] ),
    .S0(net442),
    .S1(net450),
    .X(_11133_));
 sky130_fd_sc_hd__mux4_2 _25317_ (.A0(\w[16][13] ),
    .A1(\w[20][13] ),
    .A2(\w[18][13] ),
    .A3(\w[22][13] ),
    .S0(net442),
    .S1(net450),
    .X(_11134_));
 sky130_fd_sc_hd__mux4_2 _25318_ (.A0(\w[24][13] ),
    .A1(\w[28][13] ),
    .A2(\w[26][13] ),
    .A3(\w[30][13] ),
    .S0(net442),
    .S1(net450),
    .X(_11135_));
 sky130_fd_sc_hd__mux4_2 _25319_ (.A0(_11132_),
    .A1(_11133_),
    .A2(_11134_),
    .A3(_11135_),
    .S0(net437),
    .S1(net435),
    .X(_11136_));
 sky130_fd_sc_hd__mux4_2 _25320_ (.A0(\w[32][13] ),
    .A1(\w[36][13] ),
    .A2(\w[34][13] ),
    .A3(\w[38][13] ),
    .S0(net443),
    .S1(net451),
    .X(_11137_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_295 ();
 sky130_fd_sc_hd__mux4_2 _25323_ (.A0(\w[40][13] ),
    .A1(\w[44][13] ),
    .A2(\w[42][13] ),
    .A3(\w[46][13] ),
    .S0(net443),
    .S1(net451),
    .X(_11140_));
 sky130_fd_sc_hd__mux4_2 _25324_ (.A0(\w[48][13] ),
    .A1(\w[52][13] ),
    .A2(\w[50][13] ),
    .A3(\w[54][13] ),
    .S0(net445),
    .S1(net452),
    .X(_11141_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_294 ();
 sky130_fd_sc_hd__mux4_2 _25326_ (.A0(\w[56][13] ),
    .A1(\w[60][13] ),
    .A2(\w[58][13] ),
    .A3(\w[62][13] ),
    .S0(net445),
    .S1(net452),
    .X(_11143_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_293 ();
 sky130_fd_sc_hd__mux4_2 _25328_ (.A0(_11137_),
    .A1(_11140_),
    .A2(_11141_),
    .A3(_11143_),
    .S0(net438),
    .S1(net435),
    .X(_11145_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_292 ();
 sky130_fd_sc_hd__mux2i_4 _25330_ (.A0(_11136_),
    .A1(_11145_),
    .S(net432),
    .Y(_11147_));
 sky130_fd_sc_hd__mux4_2 _25331_ (.A0(\w[0][22] ),
    .A1(\w[4][22] ),
    .A2(\w[2][22] ),
    .A3(\w[6][22] ),
    .S0(net439),
    .S1(net448),
    .X(_11148_));
 sky130_fd_sc_hd__mux4_2 _25332_ (.A0(\w[8][22] ),
    .A1(\w[12][22] ),
    .A2(\w[10][22] ),
    .A3(\w[14][22] ),
    .S0(net440),
    .S1(net448),
    .X(_11149_));
 sky130_fd_sc_hd__mux4_2 _25333_ (.A0(\w[16][22] ),
    .A1(\w[20][22] ),
    .A2(\w[18][22] ),
    .A3(\w[22][22] ),
    .S0(net440),
    .S1(net448),
    .X(_11150_));
 sky130_fd_sc_hd__mux4_2 _25334_ (.A0(\w[24][22] ),
    .A1(\w[28][22] ),
    .A2(\w[26][22] ),
    .A3(\w[30][22] ),
    .S0(net440),
    .S1(net448),
    .X(_11151_));
 sky130_fd_sc_hd__mux4_2 _25335_ (.A0(_11148_),
    .A1(_11149_),
    .A2(_11150_),
    .A3(_11151_),
    .S0(net436),
    .S1(net434),
    .X(_11152_));
 sky130_fd_sc_hd__mux4_2 _25336_ (.A0(\w[32][22] ),
    .A1(\w[36][22] ),
    .A2(\w[34][22] ),
    .A3(\w[38][22] ),
    .S0(net439),
    .S1(net448),
    .X(_11153_));
 sky130_fd_sc_hd__mux4_2 _25337_ (.A0(\w[40][22] ),
    .A1(\w[44][22] ),
    .A2(\w[42][22] ),
    .A3(\w[46][22] ),
    .S0(net439),
    .S1(net448),
    .X(_11154_));
 sky130_fd_sc_hd__mux4_2 _25338_ (.A0(\w[48][22] ),
    .A1(\w[52][22] ),
    .A2(\w[50][22] ),
    .A3(\w[54][22] ),
    .S0(net439),
    .S1(net448),
    .X(_11155_));
 sky130_fd_sc_hd__mux4_2 _25339_ (.A0(\w[56][22] ),
    .A1(\w[60][22] ),
    .A2(\w[58][22] ),
    .A3(\w[62][22] ),
    .S0(net439),
    .S1(net448),
    .X(_11156_));
 sky130_fd_sc_hd__mux4_2 _25340_ (.A0(_11153_),
    .A1(_11154_),
    .A2(_11155_),
    .A3(_11156_),
    .S0(net436),
    .S1(net434),
    .X(_11157_));
 sky130_fd_sc_hd__mux2i_4 _25341_ (.A0(_11152_),
    .A1(_11157_),
    .S(net432),
    .Y(_11158_));
 sky130_fd_sc_hd__xnor2_1 _25342_ (.A(_11147_),
    .B(_11158_),
    .Y(_11159_));
 sky130_fd_sc_hd__xnor2_1 _25343_ (.A(_10995_),
    .B(_11159_),
    .Y(_11608_));
 sky130_fd_sc_hd__mux4_2 _25344_ (.A0(\w[1][22] ),
    .A1(\w[5][22] ),
    .A2(\w[3][22] ),
    .A3(\w[7][22] ),
    .S0(net524),
    .S1(net529),
    .X(_11160_));
 sky130_fd_sc_hd__mux4_2 _25345_ (.A0(\w[9][22] ),
    .A1(\w[13][22] ),
    .A2(\w[11][22] ),
    .A3(\w[15][22] ),
    .S0(net524),
    .S1(net529),
    .X(_11161_));
 sky130_fd_sc_hd__mux4_2 _25346_ (.A0(\w[17][22] ),
    .A1(\w[21][22] ),
    .A2(\w[19][22] ),
    .A3(\w[23][22] ),
    .S0(net524),
    .S1(net529),
    .X(_11162_));
 sky130_fd_sc_hd__mux4_2 _25347_ (.A0(\w[25][22] ),
    .A1(\w[29][22] ),
    .A2(\w[27][22] ),
    .A3(\w[31][22] ),
    .S0(net524),
    .S1(net529),
    .X(_11163_));
 sky130_fd_sc_hd__mux4_2 _25348_ (.A0(_11160_),
    .A1(_11161_),
    .A2(_11162_),
    .A3(_11163_),
    .S0(net517),
    .S1(net515),
    .X(_11164_));
 sky130_fd_sc_hd__mux4_2 _25349_ (.A0(\w[33][22] ),
    .A1(\w[37][22] ),
    .A2(\w[35][22] ),
    .A3(\w[39][22] ),
    .S0(net525),
    .S1(net529),
    .X(_11165_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_291 ();
 sky130_fd_sc_hd__mux4_2 _25351_ (.A0(\w[41][22] ),
    .A1(\w[45][22] ),
    .A2(\w[43][22] ),
    .A3(\w[47][22] ),
    .S0(net525),
    .S1(net529),
    .X(_11167_));
 sky130_fd_sc_hd__mux4_2 _25352_ (.A0(\w[49][22] ),
    .A1(\w[53][22] ),
    .A2(\w[51][22] ),
    .A3(\w[55][22] ),
    .S0(net525),
    .S1(net529),
    .X(_11168_));
 sky130_fd_sc_hd__mux4_2 _25353_ (.A0(\w[57][22] ),
    .A1(\w[61][22] ),
    .A2(\w[59][22] ),
    .A3(\w[63][22] ),
    .S0(net525),
    .S1(net529),
    .X(_11169_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_290 ();
 sky130_fd_sc_hd__mux4_2 _25355_ (.A0(_11165_),
    .A1(_11167_),
    .A2(_11168_),
    .A3(_11169_),
    .S0(net517),
    .S1(net515),
    .X(_11171_));
 sky130_fd_sc_hd__mux2i_4 _25356_ (.A0(_11164_),
    .A1(_11171_),
    .S(\count15_1[5] ),
    .Y(_11172_));
 sky130_fd_sc_hd__mux4_2 _25357_ (.A0(\w[1][11] ),
    .A1(\w[5][11] ),
    .A2(\w[3][11] ),
    .A3(\w[7][11] ),
    .S0(net525),
    .S1(net529),
    .X(_11173_));
 sky130_fd_sc_hd__mux4_2 _25358_ (.A0(\w[9][11] ),
    .A1(\w[13][11] ),
    .A2(\w[11][11] ),
    .A3(\w[15][11] ),
    .S0(net525),
    .S1(net529),
    .X(_11174_));
 sky130_fd_sc_hd__mux4_2 _25359_ (.A0(\w[17][11] ),
    .A1(\w[21][11] ),
    .A2(\w[19][11] ),
    .A3(\w[23][11] ),
    .S0(net525),
    .S1(net529),
    .X(_11175_));
 sky130_fd_sc_hd__mux4_2 _25360_ (.A0(\w[25][11] ),
    .A1(\w[29][11] ),
    .A2(\w[27][11] ),
    .A3(\w[31][11] ),
    .S0(net525),
    .S1(net529),
    .X(_11176_));
 sky130_fd_sc_hd__mux4_2 _25361_ (.A0(_11173_),
    .A1(_11174_),
    .A2(_11175_),
    .A3(_11176_),
    .S0(net517),
    .S1(net514),
    .X(_11177_));
 sky130_fd_sc_hd__mux4_2 _25362_ (.A0(\w[33][11] ),
    .A1(\w[37][11] ),
    .A2(\w[35][11] ),
    .A3(\w[39][11] ),
    .S0(net527),
    .S1(net550),
    .X(_11178_));
 sky130_fd_sc_hd__mux4_2 _25363_ (.A0(\w[41][11] ),
    .A1(\w[45][11] ),
    .A2(\w[43][11] ),
    .A3(\w[47][11] ),
    .S0(net527),
    .S1(net550),
    .X(_11179_));
 sky130_fd_sc_hd__mux4_2 _25364_ (.A0(\w[49][11] ),
    .A1(\w[53][11] ),
    .A2(\w[51][11] ),
    .A3(\w[55][11] ),
    .S0(net527),
    .S1(net550),
    .X(_11180_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_289 ();
 sky130_fd_sc_hd__mux4_2 _25366_ (.A0(\w[57][11] ),
    .A1(\w[61][11] ),
    .A2(\w[59][11] ),
    .A3(\w[63][11] ),
    .S0(net527),
    .S1(net550),
    .X(_11182_));
 sky130_fd_sc_hd__mux4_2 _25367_ (.A0(_11178_),
    .A1(_11179_),
    .A2(_11180_),
    .A3(_11182_),
    .S0(\count15_1[3] ),
    .S1(net515),
    .X(_11183_));
 sky130_fd_sc_hd__mux2i_4 _25368_ (.A0(_11177_),
    .A1(_11183_),
    .S(\count15_1[5] ),
    .Y(_11184_));
 sky130_fd_sc_hd__xnor2_1 _25369_ (.A(_11172_),
    .B(_11184_),
    .Y(_11185_));
 sky130_fd_sc_hd__xnor2_1 _25370_ (.A(_10893_),
    .B(_11185_),
    .Y(_11611_));
 sky130_fd_sc_hd__mux4_2 _25371_ (.A0(\w[0][14] ),
    .A1(\w[4][14] ),
    .A2(\w[2][14] ),
    .A3(\w[6][14] ),
    .S0(net445),
    .S1(net452),
    .X(_11186_));
 sky130_fd_sc_hd__mux4_2 _25372_ (.A0(\w[8][14] ),
    .A1(\w[12][14] ),
    .A2(\w[10][14] ),
    .A3(\w[14][14] ),
    .S0(net445),
    .S1(net452),
    .X(_11187_));
 sky130_fd_sc_hd__mux4_2 _25373_ (.A0(\w[16][14] ),
    .A1(\w[20][14] ),
    .A2(\w[18][14] ),
    .A3(\w[22][14] ),
    .S0(net445),
    .S1(net452),
    .X(_11188_));
 sky130_fd_sc_hd__mux4_2 _25374_ (.A0(\w[24][14] ),
    .A1(\w[28][14] ),
    .A2(\w[26][14] ),
    .A3(\w[30][14] ),
    .S0(net445),
    .S1(net452),
    .X(_11189_));
 sky130_fd_sc_hd__mux4_2 _25375_ (.A0(_11186_),
    .A1(_11187_),
    .A2(_11188_),
    .A3(_11189_),
    .S0(net437),
    .S1(net435),
    .X(_11190_));
 sky130_fd_sc_hd__mux4_2 _25376_ (.A0(\w[32][14] ),
    .A1(\w[36][14] ),
    .A2(\w[34][14] ),
    .A3(\w[38][14] ),
    .S0(net443),
    .S1(net451),
    .X(_11191_));
 sky130_fd_sc_hd__mux4_2 _25377_ (.A0(\w[40][14] ),
    .A1(\w[44][14] ),
    .A2(\w[42][14] ),
    .A3(\w[46][14] ),
    .S0(net443),
    .S1(net451),
    .X(_11192_));
 sky130_fd_sc_hd__mux4_2 _25378_ (.A0(\w[48][14] ),
    .A1(\w[52][14] ),
    .A2(\w[50][14] ),
    .A3(\w[54][14] ),
    .S0(net443),
    .S1(net451),
    .X(_11193_));
 sky130_fd_sc_hd__mux4_2 _25379_ (.A0(\w[56][14] ),
    .A1(\w[60][14] ),
    .A2(\w[58][14] ),
    .A3(\w[62][14] ),
    .S0(net443),
    .S1(net451),
    .X(_11194_));
 sky130_fd_sc_hd__mux4_2 _25380_ (.A0(_11191_),
    .A1(_11192_),
    .A2(_11193_),
    .A3(_11194_),
    .S0(net438),
    .S1(net435),
    .X(_11195_));
 sky130_fd_sc_hd__mux2i_4 _25381_ (.A0(_11190_),
    .A1(_11195_),
    .S(net432),
    .Y(_11196_));
 sky130_fd_sc_hd__mux4_2 _25382_ (.A0(\w[0][23] ),
    .A1(\w[4][23] ),
    .A2(\w[2][23] ),
    .A3(\w[6][23] ),
    .S0(net445),
    .S1(net452),
    .X(_11197_));
 sky130_fd_sc_hd__mux4_2 _25383_ (.A0(\w[8][23] ),
    .A1(\w[12][23] ),
    .A2(\w[10][23] ),
    .A3(\w[14][23] ),
    .S0(net445),
    .S1(net452),
    .X(_11198_));
 sky130_fd_sc_hd__mux4_2 _25384_ (.A0(\w[16][23] ),
    .A1(\w[20][23] ),
    .A2(\w[18][23] ),
    .A3(\w[22][23] ),
    .S0(net445),
    .S1(net452),
    .X(_11199_));
 sky130_fd_sc_hd__mux4_2 _25385_ (.A0(\w[24][23] ),
    .A1(\w[28][23] ),
    .A2(\w[26][23] ),
    .A3(\w[30][23] ),
    .S0(net445),
    .S1(net452),
    .X(_11200_));
 sky130_fd_sc_hd__mux4_2 _25386_ (.A0(_11197_),
    .A1(_11198_),
    .A2(_11199_),
    .A3(_11200_),
    .S0(net437),
    .S1(net435),
    .X(_11201_));
 sky130_fd_sc_hd__mux4_2 _25387_ (.A0(\w[32][23] ),
    .A1(\w[36][23] ),
    .A2(\w[34][23] ),
    .A3(\w[38][23] ),
    .S0(net442),
    .S1(net450),
    .X(_11202_));
 sky130_fd_sc_hd__mux4_2 _25388_ (.A0(\w[40][23] ),
    .A1(\w[44][23] ),
    .A2(\w[42][23] ),
    .A3(\w[46][23] ),
    .S0(net442),
    .S1(net450),
    .X(_11203_));
 sky130_fd_sc_hd__mux4_2 _25389_ (.A0(\w[48][23] ),
    .A1(\w[52][23] ),
    .A2(\w[50][23] ),
    .A3(\w[54][23] ),
    .S0(net442),
    .S1(net450),
    .X(_11204_));
 sky130_fd_sc_hd__mux4_2 _25390_ (.A0(\w[56][23] ),
    .A1(\w[60][23] ),
    .A2(\w[58][23] ),
    .A3(\w[62][23] ),
    .S0(net442),
    .S1(net450),
    .X(_11205_));
 sky130_fd_sc_hd__mux4_2 _25391_ (.A0(_11202_),
    .A1(_11203_),
    .A2(_11204_),
    .A3(_11205_),
    .S0(net437),
    .S1(net435),
    .X(_11206_));
 sky130_fd_sc_hd__mux2i_4 _25392_ (.A0(_11201_),
    .A1(_11206_),
    .S(net433),
    .Y(_11207_));
 sky130_fd_sc_hd__xnor2_1 _25393_ (.A(_11196_),
    .B(_11207_),
    .Y(_11208_));
 sky130_fd_sc_hd__xnor2_1 _25394_ (.A(_11071_),
    .B(_11208_),
    .Y(_11616_));
 sky130_fd_sc_hd__mux4_2 _25395_ (.A0(\w[1][23] ),
    .A1(\w[5][23] ),
    .A2(\w[3][23] ),
    .A3(\w[7][23] ),
    .S0(net523),
    .S1(net532),
    .X(_11209_));
 sky130_fd_sc_hd__mux4_2 _25396_ (.A0(\w[9][23] ),
    .A1(\w[13][23] ),
    .A2(\w[11][23] ),
    .A3(\w[15][23] ),
    .S0(net523),
    .S1(net532),
    .X(_11210_));
 sky130_fd_sc_hd__mux4_2 _25397_ (.A0(\w[17][23] ),
    .A1(\w[21][23] ),
    .A2(\w[19][23] ),
    .A3(\w[23][23] ),
    .S0(net523),
    .S1(net532),
    .X(_11211_));
 sky130_fd_sc_hd__mux4_2 _25398_ (.A0(\w[25][23] ),
    .A1(\w[29][23] ),
    .A2(\w[27][23] ),
    .A3(\w[31][23] ),
    .S0(net523),
    .S1(net532),
    .X(_11212_));
 sky130_fd_sc_hd__mux4_2 _25399_ (.A0(_11209_),
    .A1(_11210_),
    .A2(_11211_),
    .A3(_11212_),
    .S0(net518),
    .S1(net549),
    .X(_11213_));
 sky130_fd_sc_hd__mux4_2 _25400_ (.A0(\w[33][23] ),
    .A1(\w[37][23] ),
    .A2(\w[35][23] ),
    .A3(\w[39][23] ),
    .S0(net522),
    .S1(net531),
    .X(_11214_));
 sky130_fd_sc_hd__mux4_2 _25401_ (.A0(\w[41][23] ),
    .A1(\w[45][23] ),
    .A2(\w[43][23] ),
    .A3(\w[47][23] ),
    .S0(net522),
    .S1(net531),
    .X(_11215_));
 sky130_fd_sc_hd__mux4_2 _25402_ (.A0(\w[49][23] ),
    .A1(\w[53][23] ),
    .A2(\w[51][23] ),
    .A3(\w[55][23] ),
    .S0(net522),
    .S1(net531),
    .X(_11216_));
 sky130_fd_sc_hd__mux4_2 _25403_ (.A0(\w[57][23] ),
    .A1(\w[61][23] ),
    .A2(\w[59][23] ),
    .A3(\w[63][23] ),
    .S0(net522),
    .S1(net531),
    .X(_11217_));
 sky130_fd_sc_hd__mux4_2 _25404_ (.A0(_11214_),
    .A1(_11215_),
    .A2(_11216_),
    .A3(_11217_),
    .S0(net516),
    .S1(net514),
    .X(_11218_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_288 ();
 sky130_fd_sc_hd__mux2i_4 _25406_ (.A0(_11213_),
    .A1(_11218_),
    .S(net512),
    .Y(_11220_));
 sky130_fd_sc_hd__mux4_2 _25407_ (.A0(\w[1][12] ),
    .A1(\w[5][12] ),
    .A2(\w[3][12] ),
    .A3(\w[7][12] ),
    .S0(net525),
    .S1(net529),
    .X(_11221_));
 sky130_fd_sc_hd__mux4_2 _25408_ (.A0(\w[9][12] ),
    .A1(\w[13][12] ),
    .A2(\w[11][12] ),
    .A3(\w[15][12] ),
    .S0(net525),
    .S1(net529),
    .X(_11222_));
 sky130_fd_sc_hd__mux4_2 _25409_ (.A0(\w[17][12] ),
    .A1(\w[21][12] ),
    .A2(\w[19][12] ),
    .A3(\w[23][12] ),
    .S0(net525),
    .S1(net529),
    .X(_11223_));
 sky130_fd_sc_hd__mux4_2 _25410_ (.A0(\w[25][12] ),
    .A1(\w[29][12] ),
    .A2(\w[27][12] ),
    .A3(\w[31][12] ),
    .S0(net525),
    .S1(net529),
    .X(_11224_));
 sky130_fd_sc_hd__mux4_2 _25411_ (.A0(_11221_),
    .A1(_11222_),
    .A2(_11223_),
    .A3(_11224_),
    .S0(net517),
    .S1(net515),
    .X(_11225_));
 sky130_fd_sc_hd__mux4_2 _25412_ (.A0(\w[33][12] ),
    .A1(\w[37][12] ),
    .A2(\w[35][12] ),
    .A3(\w[39][12] ),
    .S0(net526),
    .S1(net530),
    .X(_11226_));
 sky130_fd_sc_hd__mux4_2 _25413_ (.A0(\w[41][12] ),
    .A1(\w[45][12] ),
    .A2(\w[43][12] ),
    .A3(\w[47][12] ),
    .S0(net526),
    .S1(net530),
    .X(_11227_));
 sky130_fd_sc_hd__mux4_2 _25414_ (.A0(\w[49][12] ),
    .A1(\w[53][12] ),
    .A2(\w[51][12] ),
    .A3(\w[55][12] ),
    .S0(net526),
    .S1(net530),
    .X(_11228_));
 sky130_fd_sc_hd__mux4_2 _25415_ (.A0(\w[57][12] ),
    .A1(\w[61][12] ),
    .A2(\w[59][12] ),
    .A3(\w[63][12] ),
    .S0(net526),
    .S1(net530),
    .X(_11229_));
 sky130_fd_sc_hd__mux4_2 _25416_ (.A0(_11226_),
    .A1(_11227_),
    .A2(_11228_),
    .A3(_11229_),
    .S0(net517),
    .S1(net515),
    .X(_11230_));
 sky130_fd_sc_hd__mux2i_4 _25417_ (.A0(_11225_),
    .A1(_11230_),
    .S(\count15_1[5] ),
    .Y(_11231_));
 sky130_fd_sc_hd__xnor2_1 _25418_ (.A(_11220_),
    .B(_11231_),
    .Y(_11232_));
 sky130_fd_sc_hd__xnor2_1 _25419_ (.A(_10917_),
    .B(_11232_),
    .Y(_11619_));
 sky130_fd_sc_hd__mux4_2 _25420_ (.A0(\w[0][15] ),
    .A1(\w[4][15] ),
    .A2(\w[2][15] ),
    .A3(\w[6][15] ),
    .S0(net446),
    .S1(net447),
    .X(_11233_));
 sky130_fd_sc_hd__mux4_2 _25421_ (.A0(\w[8][15] ),
    .A1(\w[12][15] ),
    .A2(\w[10][15] ),
    .A3(\w[14][15] ),
    .S0(net446),
    .S1(net447),
    .X(_11234_));
 sky130_fd_sc_hd__mux4_2 _25422_ (.A0(\w[16][15] ),
    .A1(\w[20][15] ),
    .A2(\w[18][15] ),
    .A3(\w[22][15] ),
    .S0(net446),
    .S1(net447),
    .X(_11235_));
 sky130_fd_sc_hd__mux4_2 _25423_ (.A0(\w[24][15] ),
    .A1(\w[28][15] ),
    .A2(\w[26][15] ),
    .A3(\w[30][15] ),
    .S0(net446),
    .S1(net447),
    .X(_11236_));
 sky130_fd_sc_hd__mux4_2 _25424_ (.A0(_11233_),
    .A1(_11234_),
    .A2(_11235_),
    .A3(_11236_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_11237_));
 sky130_fd_sc_hd__mux4_2 _25425_ (.A0(\w[32][15] ),
    .A1(\w[36][15] ),
    .A2(\w[34][15] ),
    .A3(\w[38][15] ),
    .S0(net446),
    .S1(net1093),
    .X(_11238_));
 sky130_fd_sc_hd__mux4_2 _25426_ (.A0(\w[40][15] ),
    .A1(\w[44][15] ),
    .A2(\w[42][15] ),
    .A3(\w[46][15] ),
    .S0(net446),
    .S1(net447),
    .X(_11239_));
 sky130_fd_sc_hd__mux4_2 _25427_ (.A0(\w[48][15] ),
    .A1(\w[52][15] ),
    .A2(\w[50][15] ),
    .A3(\w[54][15] ),
    .S0(net446),
    .S1(net447),
    .X(_11240_));
 sky130_fd_sc_hd__mux4_2 _25428_ (.A0(\w[56][15] ),
    .A1(\w[60][15] ),
    .A2(\w[58][15] ),
    .A3(\w[62][15] ),
    .S0(net446),
    .S1(net447),
    .X(_11241_));
 sky130_fd_sc_hd__mux4_2 _25429_ (.A0(_11238_),
    .A1(_11239_),
    .A2(_11240_),
    .A3(_11241_),
    .S0(net437),
    .S1(net435),
    .X(_11242_));
 sky130_fd_sc_hd__mux2i_4 _25430_ (.A0(_11237_),
    .A1(_11242_),
    .S(\count2_1[5] ),
    .Y(_11243_));
 sky130_fd_sc_hd__mux4_2 _25431_ (.A0(\w[0][24] ),
    .A1(\w[4][24] ),
    .A2(\w[2][24] ),
    .A3(\w[6][24] ),
    .S0(net439),
    .S1(net448),
    .X(_11244_));
 sky130_fd_sc_hd__mux4_2 _25432_ (.A0(\w[8][24] ),
    .A1(\w[12][24] ),
    .A2(\w[10][24] ),
    .A3(\w[14][24] ),
    .S0(net439),
    .S1(net448),
    .X(_11245_));
 sky130_fd_sc_hd__mux4_2 _25433_ (.A0(\w[16][24] ),
    .A1(\w[20][24] ),
    .A2(\w[18][24] ),
    .A3(\w[22][24] ),
    .S0(net439),
    .S1(net448),
    .X(_11246_));
 sky130_fd_sc_hd__mux4_2 _25434_ (.A0(\w[24][24] ),
    .A1(\w[28][24] ),
    .A2(\w[26][24] ),
    .A3(\w[30][24] ),
    .S0(net439),
    .S1(net448),
    .X(_11247_));
 sky130_fd_sc_hd__mux4_2 _25435_ (.A0(_11244_),
    .A1(_11245_),
    .A2(_11246_),
    .A3(_11247_),
    .S0(net436),
    .S1(net434),
    .X(_11248_));
 sky130_fd_sc_hd__mux4_2 _25436_ (.A0(\w[32][24] ),
    .A1(\w[36][24] ),
    .A2(\w[34][24] ),
    .A3(\w[38][24] ),
    .S0(net440),
    .S1(net448),
    .X(_11249_));
 sky130_fd_sc_hd__mux4_2 _25437_ (.A0(\w[40][24] ),
    .A1(\w[44][24] ),
    .A2(\w[42][24] ),
    .A3(\w[46][24] ),
    .S0(net439),
    .S1(net448),
    .X(_11250_));
 sky130_fd_sc_hd__mux4_2 _25438_ (.A0(\w[48][24] ),
    .A1(\w[52][24] ),
    .A2(\w[50][24] ),
    .A3(\w[54][24] ),
    .S0(net440),
    .S1(net448),
    .X(_11251_));
 sky130_fd_sc_hd__mux4_2 _25439_ (.A0(\w[56][24] ),
    .A1(\w[60][24] ),
    .A2(\w[58][24] ),
    .A3(\w[62][24] ),
    .S0(net440),
    .S1(net448),
    .X(_11252_));
 sky130_fd_sc_hd__mux4_2 _25440_ (.A0(_11249_),
    .A1(_11250_),
    .A2(_11251_),
    .A3(_11252_),
    .S0(net438),
    .S1(net434),
    .X(_11253_));
 sky130_fd_sc_hd__mux2i_4 _25441_ (.A0(_11248_),
    .A1(_11253_),
    .S(net432),
    .Y(_11254_));
 sky130_fd_sc_hd__xnor2_1 _25442_ (.A(_11243_),
    .B(_11254_),
    .Y(_11255_));
 sky130_fd_sc_hd__xnor2_1 _25443_ (.A(_11158_),
    .B(_11255_),
    .Y(_11624_));
 sky130_fd_sc_hd__mux4_2 _25444_ (.A0(\w[1][24] ),
    .A1(\w[5][24] ),
    .A2(\w[3][24] ),
    .A3(\w[7][24] ),
    .S0(net521),
    .S1(net528),
    .X(_11256_));
 sky130_fd_sc_hd__mux4_2 _25445_ (.A0(\w[9][24] ),
    .A1(\w[13][24] ),
    .A2(\w[11][24] ),
    .A3(\w[15][24] ),
    .S0(net521),
    .S1(net528),
    .X(_11257_));
 sky130_fd_sc_hd__mux4_2 _25446_ (.A0(\w[17][24] ),
    .A1(\w[21][24] ),
    .A2(\w[19][24] ),
    .A3(\w[23][24] ),
    .S0(net521),
    .S1(net528),
    .X(_11258_));
 sky130_fd_sc_hd__mux4_2 _25447_ (.A0(\w[25][24] ),
    .A1(\w[29][24] ),
    .A2(\w[27][24] ),
    .A3(\w[31][24] ),
    .S0(net521),
    .S1(net528),
    .X(_11259_));
 sky130_fd_sc_hd__mux4_2 _25448_ (.A0(_11256_),
    .A1(_11257_),
    .A2(_11258_),
    .A3(_11259_),
    .S0(net516),
    .S1(net514),
    .X(_11260_));
 sky130_fd_sc_hd__mux4_2 _25449_ (.A0(\w[33][24] ),
    .A1(\w[37][24] ),
    .A2(\w[35][24] ),
    .A3(\w[39][24] ),
    .S0(net522),
    .S1(net531),
    .X(_11261_));
 sky130_fd_sc_hd__mux4_2 _25450_ (.A0(\w[41][24] ),
    .A1(\w[45][24] ),
    .A2(\w[43][24] ),
    .A3(\w[47][24] ),
    .S0(net522),
    .S1(net530),
    .X(_11262_));
 sky130_fd_sc_hd__mux4_2 _25451_ (.A0(\w[49][24] ),
    .A1(\w[53][24] ),
    .A2(\w[51][24] ),
    .A3(\w[55][24] ),
    .S0(net522),
    .S1(net531),
    .X(_11263_));
 sky130_fd_sc_hd__mux4_2 _25452_ (.A0(\w[57][24] ),
    .A1(\w[61][24] ),
    .A2(\w[59][24] ),
    .A3(\w[63][24] ),
    .S0(net522),
    .S1(net530),
    .X(_11264_));
 sky130_fd_sc_hd__mux4_2 _25453_ (.A0(_11261_),
    .A1(_11262_),
    .A2(_11263_),
    .A3(_11264_),
    .S0(net516),
    .S1(net514),
    .X(_11265_));
 sky130_fd_sc_hd__mux2i_4 _25454_ (.A0(_11260_),
    .A1(_11265_),
    .S(net512),
    .Y(_11266_));
 sky130_fd_sc_hd__mux4_2 _25455_ (.A0(\w[1][13] ),
    .A1(\w[5][13] ),
    .A2(\w[3][13] ),
    .A3(\w[7][13] ),
    .S0(net524),
    .S1(net530),
    .X(_11267_));
 sky130_fd_sc_hd__mux4_2 _25456_ (.A0(\w[9][13] ),
    .A1(\w[13][13] ),
    .A2(\w[11][13] ),
    .A3(\w[15][13] ),
    .S0(net524),
    .S1(net530),
    .X(_11268_));
 sky130_fd_sc_hd__mux4_2 _25457_ (.A0(\w[17][13] ),
    .A1(\w[21][13] ),
    .A2(\w[19][13] ),
    .A3(\w[23][13] ),
    .S0(net524),
    .S1(net530),
    .X(_11269_));
 sky130_fd_sc_hd__mux4_2 _25458_ (.A0(\w[25][13] ),
    .A1(\w[29][13] ),
    .A2(\w[27][13] ),
    .A3(\w[31][13] ),
    .S0(net524),
    .S1(net530),
    .X(_11270_));
 sky130_fd_sc_hd__mux4_2 _25459_ (.A0(_11267_),
    .A1(_11268_),
    .A2(_11269_),
    .A3(_11270_),
    .S0(net517),
    .S1(net515),
    .X(_11271_));
 sky130_fd_sc_hd__mux4_2 _25460_ (.A0(\w[33][13] ),
    .A1(\w[37][13] ),
    .A2(\w[35][13] ),
    .A3(\w[39][13] ),
    .S0(net527),
    .S1(net550),
    .X(_11272_));
 sky130_fd_sc_hd__mux4_2 _25461_ (.A0(\w[41][13] ),
    .A1(\w[45][13] ),
    .A2(\w[43][13] ),
    .A3(\w[47][13] ),
    .S0(net527),
    .S1(net550),
    .X(_11273_));
 sky130_fd_sc_hd__mux4_2 _25462_ (.A0(\w[49][13] ),
    .A1(\w[53][13] ),
    .A2(\w[51][13] ),
    .A3(\w[55][13] ),
    .S0(net527),
    .S1(net550),
    .X(_11274_));
 sky130_fd_sc_hd__mux4_2 _25463_ (.A0(\w[57][13] ),
    .A1(\w[61][13] ),
    .A2(\w[59][13] ),
    .A3(\w[63][13] ),
    .S0(net527),
    .S1(net550),
    .X(_11275_));
 sky130_fd_sc_hd__mux4_2 _25464_ (.A0(_11272_),
    .A1(_11273_),
    .A2(_11274_),
    .A3(_11275_),
    .S0(\count15_1[3] ),
    .S1(net515),
    .X(_11276_));
 sky130_fd_sc_hd__mux2i_4 _25465_ (.A0(_11271_),
    .A1(_11276_),
    .S(\count15_1[5] ),
    .Y(_11277_));
 sky130_fd_sc_hd__xnor2_1 _25466_ (.A(_11266_),
    .B(_11277_),
    .Y(_11278_));
 sky130_fd_sc_hd__xnor2_1 _25467_ (.A(_11045_),
    .B(_11278_),
    .Y(_11627_));
 sky130_fd_sc_hd__mux4_2 _25468_ (.A0(\w[0][25] ),
    .A1(\w[4][25] ),
    .A2(\w[2][25] ),
    .A3(\w[6][25] ),
    .S0(net442),
    .S1(net450),
    .X(_11279_));
 sky130_fd_sc_hd__mux4_2 _25469_ (.A0(\w[8][25] ),
    .A1(\w[12][25] ),
    .A2(\w[10][25] ),
    .A3(\w[14][25] ),
    .S0(net442),
    .S1(net450),
    .X(_11280_));
 sky130_fd_sc_hd__mux4_2 _25470_ (.A0(\w[16][25] ),
    .A1(\w[20][25] ),
    .A2(\w[18][25] ),
    .A3(\w[22][25] ),
    .S0(net442),
    .S1(net450),
    .X(_11281_));
 sky130_fd_sc_hd__mux4_2 _25471_ (.A0(\w[24][25] ),
    .A1(\w[28][25] ),
    .A2(\w[26][25] ),
    .A3(\w[30][25] ),
    .S0(net442),
    .S1(net450),
    .X(_11282_));
 sky130_fd_sc_hd__mux4_2 _25472_ (.A0(_11279_),
    .A1(_11280_),
    .A2(_11281_),
    .A3(_11282_),
    .S0(net438),
    .S1(net434),
    .X(_11283_));
 sky130_fd_sc_hd__mux4_2 _25473_ (.A0(\w[32][25] ),
    .A1(\w[36][25] ),
    .A2(\w[34][25] ),
    .A3(\w[38][25] ),
    .S0(net441),
    .S1(net449),
    .X(_11284_));
 sky130_fd_sc_hd__mux4_2 _25474_ (.A0(\w[40][25] ),
    .A1(\w[44][25] ),
    .A2(\w[42][25] ),
    .A3(\w[46][25] ),
    .S0(net441),
    .S1(net449),
    .X(_11285_));
 sky130_fd_sc_hd__mux4_2 _25475_ (.A0(\w[48][25] ),
    .A1(\w[52][25] ),
    .A2(\w[50][25] ),
    .A3(\w[54][25] ),
    .S0(net441),
    .S1(net449),
    .X(_11286_));
 sky130_fd_sc_hd__mux4_2 _25476_ (.A0(\w[56][25] ),
    .A1(\w[60][25] ),
    .A2(\w[58][25] ),
    .A3(\w[62][25] ),
    .S0(net441),
    .S1(net449),
    .X(_11287_));
 sky130_fd_sc_hd__mux4_2 _25477_ (.A0(_11284_),
    .A1(_11285_),
    .A2(_11286_),
    .A3(_11287_),
    .S0(net438),
    .S1(net434),
    .X(_11288_));
 sky130_fd_sc_hd__mux2i_4 _25478_ (.A0(_11283_),
    .A1(_11288_),
    .S(net432),
    .Y(_11289_));
 sky130_fd_sc_hd__mux4_2 _25479_ (.A0(\w[0][16] ),
    .A1(\w[4][16] ),
    .A2(\w[2][16] ),
    .A3(\w[6][16] ),
    .S0(net446),
    .S1(net447),
    .X(_11290_));
 sky130_fd_sc_hd__mux4_2 _25480_ (.A0(\w[8][16] ),
    .A1(\w[12][16] ),
    .A2(\w[10][16] ),
    .A3(\w[14][16] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_11291_));
 sky130_fd_sc_hd__mux4_2 _25481_ (.A0(\w[16][16] ),
    .A1(\w[20][16] ),
    .A2(\w[18][16] ),
    .A3(\w[22][16] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_11292_));
 sky130_fd_sc_hd__mux4_2 _25482_ (.A0(\w[24][16] ),
    .A1(\w[28][16] ),
    .A2(\w[26][16] ),
    .A3(\w[30][16] ),
    .S0(net446),
    .S1(net447),
    .X(_11293_));
 sky130_fd_sc_hd__mux4_2 _25483_ (.A0(_11290_),
    .A1(_11291_),
    .A2(_11292_),
    .A3(_11293_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_11294_));
 sky130_fd_sc_hd__mux4_2 _25484_ (.A0(\w[32][16] ),
    .A1(\w[36][16] ),
    .A2(\w[34][16] ),
    .A3(\w[38][16] ),
    .S0(\count2_1[2] ),
    .S1(net452),
    .X(_11295_));
 sky130_fd_sc_hd__mux4_2 _25485_ (.A0(\w[40][16] ),
    .A1(\w[44][16] ),
    .A2(\w[42][16] ),
    .A3(\w[46][16] ),
    .S0(\count2_1[2] ),
    .S1(net452),
    .X(_11296_));
 sky130_fd_sc_hd__mux4_2 _25486_ (.A0(\w[48][16] ),
    .A1(\w[52][16] ),
    .A2(\w[50][16] ),
    .A3(\w[54][16] ),
    .S0(\count2_1[2] ),
    .S1(net452),
    .X(_11297_));
 sky130_fd_sc_hd__mux4_2 _25487_ (.A0(\w[56][16] ),
    .A1(\w[60][16] ),
    .A2(\w[58][16] ),
    .A3(\w[62][16] ),
    .S0(\count2_1[2] ),
    .S1(net452),
    .X(_11298_));
 sky130_fd_sc_hd__mux4_2 _25488_ (.A0(_11295_),
    .A1(_11296_),
    .A2(_11297_),
    .A3(_11298_),
    .S0(net438),
    .S1(\count2_1[4] ),
    .X(_11299_));
 sky130_fd_sc_hd__mux2i_4 _25489_ (.A0(_11294_),
    .A1(_11299_),
    .S(net433),
    .Y(_11300_));
 sky130_fd_sc_hd__xnor2_1 _25490_ (.A(_11289_),
    .B(_11300_),
    .Y(_11301_));
 sky130_fd_sc_hd__xnor2_1 _25491_ (.A(_11207_),
    .B(_11301_),
    .Y(_11632_));
 sky130_fd_sc_hd__mux4_2 _25492_ (.A0(\w[1][14] ),
    .A1(\w[5][14] ),
    .A2(\w[3][14] ),
    .A3(\w[7][14] ),
    .S0(net526),
    .S1(net531),
    .X(_11302_));
 sky130_fd_sc_hd__mux4_2 _25493_ (.A0(\w[9][14] ),
    .A1(\w[13][14] ),
    .A2(\w[11][14] ),
    .A3(\w[15][14] ),
    .S0(net526),
    .S1(net531),
    .X(_11303_));
 sky130_fd_sc_hd__mux4_2 _25494_ (.A0(\w[17][14] ),
    .A1(\w[21][14] ),
    .A2(\w[19][14] ),
    .A3(\w[23][14] ),
    .S0(net526),
    .S1(net531),
    .X(_11304_));
 sky130_fd_sc_hd__mux4_2 _25495_ (.A0(\w[25][14] ),
    .A1(\w[29][14] ),
    .A2(\w[27][14] ),
    .A3(\w[31][14] ),
    .S0(net526),
    .S1(net531),
    .X(_11305_));
 sky130_fd_sc_hd__mux4_2 _25496_ (.A0(_11302_),
    .A1(_11303_),
    .A2(_11304_),
    .A3(_11305_),
    .S0(net517),
    .S1(net514),
    .X(_11306_));
 sky130_fd_sc_hd__mux4_2 _25497_ (.A0(\w[33][14] ),
    .A1(\w[37][14] ),
    .A2(\w[35][14] ),
    .A3(\w[39][14] ),
    .S0(net526),
    .S1(net529),
    .X(_11307_));
 sky130_fd_sc_hd__mux4_2 _25498_ (.A0(\w[41][14] ),
    .A1(\w[45][14] ),
    .A2(\w[43][14] ),
    .A3(\w[47][14] ),
    .S0(net526),
    .S1(net529),
    .X(_11308_));
 sky130_fd_sc_hd__mux4_2 _25499_ (.A0(\w[49][14] ),
    .A1(\w[53][14] ),
    .A2(\w[51][14] ),
    .A3(\w[55][14] ),
    .S0(net526),
    .S1(net529),
    .X(_11309_));
 sky130_fd_sc_hd__mux4_2 _25500_ (.A0(\w[57][14] ),
    .A1(\w[61][14] ),
    .A2(\w[59][14] ),
    .A3(\w[63][14] ),
    .S0(net526),
    .S1(net529),
    .X(_11310_));
 sky130_fd_sc_hd__mux4_2 _25501_ (.A0(_11307_),
    .A1(_11308_),
    .A2(_11309_),
    .A3(_11310_),
    .S0(net517),
    .S1(net514),
    .X(_11311_));
 sky130_fd_sc_hd__mux2i_4 _25502_ (.A0(_11306_),
    .A1(_11311_),
    .S(net512),
    .Y(_11312_));
 sky130_fd_sc_hd__mux4_2 _25503_ (.A0(\w[1][25] ),
    .A1(\w[5][25] ),
    .A2(\w[3][25] ),
    .A3(\w[7][25] ),
    .S0(net525),
    .S1(net529),
    .X(_11313_));
 sky130_fd_sc_hd__mux4_2 _25504_ (.A0(\w[9][25] ),
    .A1(\w[13][25] ),
    .A2(\w[11][25] ),
    .A3(\w[15][25] ),
    .S0(net525),
    .S1(net529),
    .X(_11314_));
 sky130_fd_sc_hd__mux4_2 _25505_ (.A0(\w[17][25] ),
    .A1(\w[21][25] ),
    .A2(\w[19][25] ),
    .A3(\w[23][25] ),
    .S0(net525),
    .S1(net529),
    .X(_11315_));
 sky130_fd_sc_hd__mux4_2 _25506_ (.A0(\w[25][25] ),
    .A1(\w[29][25] ),
    .A2(\w[27][25] ),
    .A3(\w[31][25] ),
    .S0(net525),
    .S1(net529),
    .X(_11316_));
 sky130_fd_sc_hd__mux4_2 _25507_ (.A0(_11313_),
    .A1(_11314_),
    .A2(_11315_),
    .A3(_11316_),
    .S0(net517),
    .S1(net515),
    .X(_11317_));
 sky130_fd_sc_hd__mux4_2 _25508_ (.A0(\w[33][25] ),
    .A1(\w[37][25] ),
    .A2(\w[35][25] ),
    .A3(\w[39][25] ),
    .S0(net526),
    .S1(net529),
    .X(_11318_));
 sky130_fd_sc_hd__mux4_2 _25509_ (.A0(\w[41][25] ),
    .A1(\w[45][25] ),
    .A2(\w[43][25] ),
    .A3(\w[47][25] ),
    .S0(net526),
    .S1(net529),
    .X(_11319_));
 sky130_fd_sc_hd__mux4_2 _25510_ (.A0(\w[49][25] ),
    .A1(\w[53][25] ),
    .A2(\w[51][25] ),
    .A3(\w[55][25] ),
    .S0(net526),
    .S1(net529),
    .X(_11320_));
 sky130_fd_sc_hd__mux4_2 _25511_ (.A0(\w[57][25] ),
    .A1(\w[61][25] ),
    .A2(\w[59][25] ),
    .A3(\w[63][25] ),
    .S0(net526),
    .S1(net529),
    .X(_11321_));
 sky130_fd_sc_hd__mux4_2 _25512_ (.A0(_11318_),
    .A1(_11319_),
    .A2(_11320_),
    .A3(_11321_),
    .S0(net517),
    .S1(net514),
    .X(_11322_));
 sky130_fd_sc_hd__mux2i_4 _25513_ (.A0(_11317_),
    .A1(_11322_),
    .S(net512),
    .Y(_11323_));
 sky130_fd_sc_hd__xnor2_1 _25514_ (.A(_11312_),
    .B(_11323_),
    .Y(_11324_));
 sky130_fd_sc_hd__xnor2_1 _25515_ (.A(_11129_),
    .B(_11324_),
    .Y(_11635_));
 sky130_fd_sc_hd__mux4_2 _25516_ (.A0(\w[0][17] ),
    .A1(\w[4][17] ),
    .A2(\w[2][17] ),
    .A3(\w[6][17] ),
    .S0(net442),
    .S1(net450),
    .X(_11325_));
 sky130_fd_sc_hd__mux4_2 _25517_ (.A0(\w[8][17] ),
    .A1(\w[12][17] ),
    .A2(\w[10][17] ),
    .A3(\w[14][17] ),
    .S0(net442),
    .S1(net450),
    .X(_11326_));
 sky130_fd_sc_hd__mux4_2 _25518_ (.A0(\w[16][17] ),
    .A1(\w[20][17] ),
    .A2(\w[18][17] ),
    .A3(\w[22][17] ),
    .S0(net442),
    .S1(net450),
    .X(_11327_));
 sky130_fd_sc_hd__mux4_2 _25519_ (.A0(\w[24][17] ),
    .A1(\w[28][17] ),
    .A2(\w[26][17] ),
    .A3(\w[30][17] ),
    .S0(net442),
    .S1(net450),
    .X(_11328_));
 sky130_fd_sc_hd__mux4_2 _25520_ (.A0(_11325_),
    .A1(_11326_),
    .A2(_11327_),
    .A3(_11328_),
    .S0(net437),
    .S1(net435),
    .X(_11329_));
 sky130_fd_sc_hd__mux4_2 _25521_ (.A0(\w[32][17] ),
    .A1(\w[36][17] ),
    .A2(\w[34][17] ),
    .A3(\w[38][17] ),
    .S0(net442),
    .S1(net450),
    .X(_11330_));
 sky130_fd_sc_hd__mux4_2 _25522_ (.A0(\w[40][17] ),
    .A1(\w[44][17] ),
    .A2(\w[42][17] ),
    .A3(\w[46][17] ),
    .S0(net442),
    .S1(net450),
    .X(_11331_));
 sky130_fd_sc_hd__mux4_2 _25523_ (.A0(\w[48][17] ),
    .A1(\w[52][17] ),
    .A2(\w[50][17] ),
    .A3(\w[54][17] ),
    .S0(net442),
    .S1(net450),
    .X(_11332_));
 sky130_fd_sc_hd__mux4_2 _25524_ (.A0(\w[56][17] ),
    .A1(\w[60][17] ),
    .A2(\w[58][17] ),
    .A3(\w[62][17] ),
    .S0(net442),
    .S1(net450),
    .X(_11333_));
 sky130_fd_sc_hd__mux4_2 _25525_ (.A0(_11330_),
    .A1(_11331_),
    .A2(_11332_),
    .A3(_11333_),
    .S0(net437),
    .S1(net435),
    .X(_11334_));
 sky130_fd_sc_hd__mux2i_4 _25526_ (.A0(_11329_),
    .A1(_11334_),
    .S(net433),
    .Y(_11335_));
 sky130_fd_sc_hd__mux4_2 _25527_ (.A0(\w[0][26] ),
    .A1(\w[4][26] ),
    .A2(\w[2][26] ),
    .A3(\w[6][26] ),
    .S0(net442),
    .S1(net450),
    .X(_11336_));
 sky130_fd_sc_hd__mux4_2 _25528_ (.A0(\w[8][26] ),
    .A1(\w[12][26] ),
    .A2(\w[10][26] ),
    .A3(\w[14][26] ),
    .S0(net442),
    .S1(net450),
    .X(_11337_));
 sky130_fd_sc_hd__mux4_2 _25529_ (.A0(\w[16][26] ),
    .A1(\w[20][26] ),
    .A2(\w[18][26] ),
    .A3(\w[22][26] ),
    .S0(net442),
    .S1(net450),
    .X(_11338_));
 sky130_fd_sc_hd__mux4_2 _25530_ (.A0(\w[24][26] ),
    .A1(\w[28][26] ),
    .A2(\w[26][26] ),
    .A3(\w[30][26] ),
    .S0(net442),
    .S1(net450),
    .X(_11339_));
 sky130_fd_sc_hd__mux4_2 _25531_ (.A0(_11336_),
    .A1(_11337_),
    .A2(_11338_),
    .A3(_11339_),
    .S0(net438),
    .S1(net434),
    .X(_11340_));
 sky130_fd_sc_hd__mux4_2 _25532_ (.A0(\w[32][26] ),
    .A1(\w[36][26] ),
    .A2(\w[34][26] ),
    .A3(\w[38][26] ),
    .S0(net441),
    .S1(net449),
    .X(_11341_));
 sky130_fd_sc_hd__mux4_2 _25533_ (.A0(\w[40][26] ),
    .A1(\w[44][26] ),
    .A2(\w[42][26] ),
    .A3(\w[46][26] ),
    .S0(net441),
    .S1(net449),
    .X(_11342_));
 sky130_fd_sc_hd__mux4_2 _25534_ (.A0(\w[48][26] ),
    .A1(\w[52][26] ),
    .A2(\w[50][26] ),
    .A3(\w[54][26] ),
    .S0(net441),
    .S1(net449),
    .X(_11343_));
 sky130_fd_sc_hd__mux4_2 _25535_ (.A0(\w[56][26] ),
    .A1(\w[60][26] ),
    .A2(\w[58][26] ),
    .A3(\w[62][26] ),
    .S0(net441),
    .S1(net449),
    .X(_11344_));
 sky130_fd_sc_hd__mux4_2 _25536_ (.A0(_11341_),
    .A1(_11342_),
    .A2(_11343_),
    .A3(_11344_),
    .S0(net438),
    .S1(net434),
    .X(_11345_));
 sky130_fd_sc_hd__mux2i_4 _25537_ (.A0(_11340_),
    .A1(_11345_),
    .S(net433),
    .Y(_11346_));
 sky130_fd_sc_hd__xnor2_1 _25538_ (.A(_11335_),
    .B(_11346_),
    .Y(_11347_));
 sky130_fd_sc_hd__xnor2_1 _25539_ (.A(_11254_),
    .B(_11347_),
    .Y(_11640_));
 sky130_fd_sc_hd__mux4_2 _25540_ (.A0(\w[1][26] ),
    .A1(\w[5][26] ),
    .A2(\w[3][26] ),
    .A3(\w[7][26] ),
    .S0(net523),
    .S1(net532),
    .X(_11348_));
 sky130_fd_sc_hd__mux4_2 _25541_ (.A0(\w[9][26] ),
    .A1(\w[13][26] ),
    .A2(\w[11][26] ),
    .A3(\w[15][26] ),
    .S0(net523),
    .S1(net532),
    .X(_11349_));
 sky130_fd_sc_hd__mux4_2 _25542_ (.A0(\w[17][26] ),
    .A1(\w[21][26] ),
    .A2(\w[19][26] ),
    .A3(\w[23][26] ),
    .S0(net523),
    .S1(net532),
    .X(_11350_));
 sky130_fd_sc_hd__mux4_2 _25543_ (.A0(\w[25][26] ),
    .A1(\w[29][26] ),
    .A2(\w[27][26] ),
    .A3(\w[31][26] ),
    .S0(net523),
    .S1(net532),
    .X(_11351_));
 sky130_fd_sc_hd__mux4_2 _25544_ (.A0(_11348_),
    .A1(_11349_),
    .A2(_11350_),
    .A3(_11351_),
    .S0(net518),
    .S1(net549),
    .X(_11352_));
 sky130_fd_sc_hd__mux4_2 _25545_ (.A0(\w[33][26] ),
    .A1(\w[37][26] ),
    .A2(\w[35][26] ),
    .A3(\w[39][26] ),
    .S0(net519),
    .S1(net531),
    .X(_11353_));
 sky130_fd_sc_hd__mux4_2 _25546_ (.A0(\w[41][26] ),
    .A1(\w[45][26] ),
    .A2(\w[43][26] ),
    .A3(\w[47][26] ),
    .S0(net519),
    .S1(net532),
    .X(_11354_));
 sky130_fd_sc_hd__mux4_2 _25547_ (.A0(\w[49][26] ),
    .A1(\w[53][26] ),
    .A2(\w[51][26] ),
    .A3(\w[55][26] ),
    .S0(net523),
    .S1(net532),
    .X(_11355_));
 sky130_fd_sc_hd__mux4_2 _25548_ (.A0(\w[57][26] ),
    .A1(\w[61][26] ),
    .A2(\w[59][26] ),
    .A3(\w[63][26] ),
    .S0(net519),
    .S1(net532),
    .X(_11356_));
 sky130_fd_sc_hd__mux4_2 _25549_ (.A0(_11353_),
    .A1(_11354_),
    .A2(_11355_),
    .A3(_11356_),
    .S0(net518),
    .S1(net549),
    .X(_11357_));
 sky130_fd_sc_hd__mux2i_4 _25550_ (.A0(_11352_),
    .A1(_11357_),
    .S(net513),
    .Y(_11358_));
 sky130_fd_sc_hd__mux4_2 _25551_ (.A0(\w[1][15] ),
    .A1(\w[5][15] ),
    .A2(\w[3][15] ),
    .A3(\w[7][15] ),
    .S0(\count15_1[2] ),
    .S1(net532),
    .X(_11359_));
 sky130_fd_sc_hd__mux4_2 _25552_ (.A0(\w[9][15] ),
    .A1(\w[13][15] ),
    .A2(\w[11][15] ),
    .A3(\w[15][15] ),
    .S0(\count15_1[2] ),
    .S1(net532),
    .X(_11360_));
 sky130_fd_sc_hd__mux4_2 _25553_ (.A0(\w[17][15] ),
    .A1(\w[21][15] ),
    .A2(\w[19][15] ),
    .A3(\w[23][15] ),
    .S0(\count15_1[2] ),
    .S1(net532),
    .X(_11361_));
 sky130_fd_sc_hd__mux4_2 _25554_ (.A0(\w[25][15] ),
    .A1(\w[29][15] ),
    .A2(\w[27][15] ),
    .A3(\w[31][15] ),
    .S0(\count15_1[2] ),
    .S1(net532),
    .X(_11362_));
 sky130_fd_sc_hd__mux4_2 _25555_ (.A0(_11359_),
    .A1(_11360_),
    .A2(_11361_),
    .A3(_11362_),
    .S0(net518),
    .S1(net549),
    .X(_11363_));
 sky130_fd_sc_hd__mux4_2 _25556_ (.A0(\w[33][15] ),
    .A1(\w[37][15] ),
    .A2(\w[35][15] ),
    .A3(\w[39][15] ),
    .S0(\count15_1[2] ),
    .S1(\count15_1[1] ),
    .X(_11364_));
 sky130_fd_sc_hd__mux4_2 _25557_ (.A0(\w[41][15] ),
    .A1(\w[45][15] ),
    .A2(\w[43][15] ),
    .A3(\w[47][15] ),
    .S0(\count15_1[2] ),
    .S1(\count15_1[1] ),
    .X(_11365_));
 sky130_fd_sc_hd__mux4_2 _25558_ (.A0(\w[49][15] ),
    .A1(\w[53][15] ),
    .A2(\w[51][15] ),
    .A3(\w[55][15] ),
    .S0(\count15_1[2] ),
    .S1(\count15_1[1] ),
    .X(_11366_));
 sky130_fd_sc_hd__mux4_2 _25559_ (.A0(\w[57][15] ),
    .A1(\w[61][15] ),
    .A2(\w[59][15] ),
    .A3(\w[63][15] ),
    .S0(\count15_1[2] ),
    .S1(\count15_1[1] ),
    .X(_11367_));
 sky130_fd_sc_hd__mux4_2 _25560_ (.A0(_11364_),
    .A1(_11365_),
    .A2(_11366_),
    .A3(_11367_),
    .S0(net518),
    .S1(net549),
    .X(_11368_));
 sky130_fd_sc_hd__mux2i_4 _25561_ (.A0(_11363_),
    .A1(_11368_),
    .S(net513),
    .Y(_11369_));
 sky130_fd_sc_hd__xnor2_1 _25562_ (.A(_11358_),
    .B(_11369_),
    .Y(_11370_));
 sky130_fd_sc_hd__xnor2_1 _25563_ (.A(_11184_),
    .B(_11370_),
    .Y(_11643_));
 sky130_fd_sc_hd__mux4_2 _25564_ (.A0(\w[0][27] ),
    .A1(\w[4][27] ),
    .A2(\w[2][27] ),
    .A3(\w[6][27] ),
    .S0(net445),
    .S1(net452),
    .X(_11371_));
 sky130_fd_sc_hd__mux4_2 _25565_ (.A0(\w[8][27] ),
    .A1(\w[12][27] ),
    .A2(\w[10][27] ),
    .A3(\w[14][27] ),
    .S0(net445),
    .S1(net452),
    .X(_11372_));
 sky130_fd_sc_hd__mux4_2 _25566_ (.A0(\w[16][27] ),
    .A1(\w[20][27] ),
    .A2(\w[18][27] ),
    .A3(\w[22][27] ),
    .S0(net445),
    .S1(net452),
    .X(_11373_));
 sky130_fd_sc_hd__mux4_2 _25567_ (.A0(\w[24][27] ),
    .A1(\w[28][27] ),
    .A2(\w[26][27] ),
    .A3(\w[30][27] ),
    .S0(net445),
    .S1(net452),
    .X(_11374_));
 sky130_fd_sc_hd__mux4_2 _25568_ (.A0(_11371_),
    .A1(_11372_),
    .A2(_11373_),
    .A3(_11374_),
    .S0(net437),
    .S1(net435),
    .X(_11375_));
 sky130_fd_sc_hd__mux4_2 _25569_ (.A0(\w[32][27] ),
    .A1(\w[36][27] ),
    .A2(\w[34][27] ),
    .A3(\w[38][27] ),
    .S0(net445),
    .S1(net452),
    .X(_11376_));
 sky130_fd_sc_hd__mux4_2 _25570_ (.A0(\w[40][27] ),
    .A1(\w[44][27] ),
    .A2(\w[42][27] ),
    .A3(\w[46][27] ),
    .S0(net445),
    .S1(net452),
    .X(_11377_));
 sky130_fd_sc_hd__mux4_2 _25571_ (.A0(\w[48][27] ),
    .A1(\w[52][27] ),
    .A2(\w[50][27] ),
    .A3(\w[54][27] ),
    .S0(net445),
    .S1(net452),
    .X(_11378_));
 sky130_fd_sc_hd__mux4_2 _25572_ (.A0(\w[56][27] ),
    .A1(\w[60][27] ),
    .A2(\w[58][27] ),
    .A3(\w[62][27] ),
    .S0(net445),
    .S1(net452),
    .X(_11379_));
 sky130_fd_sc_hd__mux4_2 _25573_ (.A0(_11376_),
    .A1(_11377_),
    .A2(_11378_),
    .A3(_11379_),
    .S0(net437),
    .S1(net435),
    .X(_11380_));
 sky130_fd_sc_hd__mux2i_4 _25574_ (.A0(_11375_),
    .A1(_11380_),
    .S(net433),
    .Y(_11381_));
 sky130_fd_sc_hd__xnor2_1 _25575_ (.A(_11289_),
    .B(_11381_),
    .Y(_11382_));
 sky130_fd_sc_hd__xnor2_1 _25576_ (.A(_11006_),
    .B(_11382_),
    .Y(_11648_));
 sky130_fd_sc_hd__mux4_2 _25577_ (.A0(\w[1][27] ),
    .A1(\w[5][27] ),
    .A2(\w[3][27] ),
    .A3(\w[7][27] ),
    .S0(net520),
    .S1(net528),
    .X(_11383_));
 sky130_fd_sc_hd__mux4_2 _25578_ (.A0(\w[9][27] ),
    .A1(\w[13][27] ),
    .A2(\w[11][27] ),
    .A3(\w[15][27] ),
    .S0(net520),
    .S1(net528),
    .X(_11384_));
 sky130_fd_sc_hd__mux4_2 _25579_ (.A0(\w[17][27] ),
    .A1(\w[21][27] ),
    .A2(\w[19][27] ),
    .A3(\w[23][27] ),
    .S0(net520),
    .S1(net528),
    .X(_11385_));
 sky130_fd_sc_hd__mux4_2 _25580_ (.A0(\w[25][27] ),
    .A1(\w[29][27] ),
    .A2(\w[27][27] ),
    .A3(\w[31][27] ),
    .S0(net520),
    .S1(net528),
    .X(_11386_));
 sky130_fd_sc_hd__mux4_2 _25581_ (.A0(_11383_),
    .A1(_11384_),
    .A2(_11385_),
    .A3(_11386_),
    .S0(net516),
    .S1(net514),
    .X(_11387_));
 sky130_fd_sc_hd__mux4_2 _25582_ (.A0(\w[33][27] ),
    .A1(\w[37][27] ),
    .A2(\w[35][27] ),
    .A3(\w[39][27] ),
    .S0(net521),
    .S1(net531),
    .X(_11388_));
 sky130_fd_sc_hd__mux4_2 _25583_ (.A0(\w[41][27] ),
    .A1(\w[45][27] ),
    .A2(\w[43][27] ),
    .A3(\w[47][27] ),
    .S0(net521),
    .S1(net531),
    .X(_11389_));
 sky130_fd_sc_hd__mux4_2 _25584_ (.A0(\w[49][27] ),
    .A1(\w[53][27] ),
    .A2(\w[51][27] ),
    .A3(\w[55][27] ),
    .S0(net521),
    .S1(net531),
    .X(_11390_));
 sky130_fd_sc_hd__mux4_2 _25585_ (.A0(\w[57][27] ),
    .A1(\w[61][27] ),
    .A2(\w[59][27] ),
    .A3(\w[63][27] ),
    .S0(net521),
    .S1(net531),
    .X(_11391_));
 sky130_fd_sc_hd__mux4_2 _25586_ (.A0(_11388_),
    .A1(_11389_),
    .A2(_11390_),
    .A3(_11391_),
    .S0(net516),
    .S1(net514),
    .X(_11392_));
 sky130_fd_sc_hd__mux2i_4 _25587_ (.A0(_11387_),
    .A1(_11392_),
    .S(net512),
    .Y(_11393_));
 sky130_fd_sc_hd__mux4_2 _25588_ (.A0(\w[1][16] ),
    .A1(\w[5][16] ),
    .A2(\w[3][16] ),
    .A3(\w[7][16] ),
    .S0(net526),
    .S1(net531),
    .X(_11394_));
 sky130_fd_sc_hd__mux4_2 _25589_ (.A0(\w[9][16] ),
    .A1(\w[13][16] ),
    .A2(\w[11][16] ),
    .A3(\w[15][16] ),
    .S0(net526),
    .S1(net531),
    .X(_11395_));
 sky130_fd_sc_hd__mux4_2 _25590_ (.A0(\w[17][16] ),
    .A1(\w[21][16] ),
    .A2(\w[19][16] ),
    .A3(\w[23][16] ),
    .S0(net522),
    .S1(net531),
    .X(_11396_));
 sky130_fd_sc_hd__mux4_2 _25591_ (.A0(\w[25][16] ),
    .A1(\w[29][16] ),
    .A2(\w[27][16] ),
    .A3(\w[31][16] ),
    .S0(net522),
    .S1(net531),
    .X(_11397_));
 sky130_fd_sc_hd__mux4_2 _25592_ (.A0(_11394_),
    .A1(_11395_),
    .A2(_11396_),
    .A3(_11397_),
    .S0(net517),
    .S1(net514),
    .X(_11398_));
 sky130_fd_sc_hd__mux4_2 _25593_ (.A0(\w[33][16] ),
    .A1(\w[37][16] ),
    .A2(\w[35][16] ),
    .A3(\w[39][16] ),
    .S0(net526),
    .S1(net530),
    .X(_11399_));
 sky130_fd_sc_hd__mux4_2 _25594_ (.A0(\w[41][16] ),
    .A1(\w[45][16] ),
    .A2(\w[43][16] ),
    .A3(\w[47][16] ),
    .S0(net526),
    .S1(net530),
    .X(_11400_));
 sky130_fd_sc_hd__mux4_2 _25595_ (.A0(\w[49][16] ),
    .A1(\w[53][16] ),
    .A2(\w[51][16] ),
    .A3(\w[55][16] ),
    .S0(net526),
    .S1(net530),
    .X(_11401_));
 sky130_fd_sc_hd__mux4_2 _25596_ (.A0(\w[57][16] ),
    .A1(\w[61][16] ),
    .A2(\w[59][16] ),
    .A3(\w[63][16] ),
    .S0(net526),
    .S1(net530),
    .X(_11402_));
 sky130_fd_sc_hd__mux4_2 _25597_ (.A0(_11399_),
    .A1(_11400_),
    .A2(_11401_),
    .A3(_11402_),
    .S0(net517),
    .S1(net514),
    .X(_11403_));
 sky130_fd_sc_hd__mux2i_4 _25598_ (.A0(_11398_),
    .A1(_11403_),
    .S(net512),
    .Y(_11404_));
 sky130_fd_sc_hd__xnor2_1 _25599_ (.A(_11393_),
    .B(_11404_),
    .Y(_11405_));
 sky130_fd_sc_hd__xnor2_1 _25600_ (.A(_11231_),
    .B(_11405_),
    .Y(_11651_));
 sky130_fd_sc_hd__mux4_2 _25601_ (.A0(\w[0][28] ),
    .A1(\w[4][28] ),
    .A2(\w[2][28] ),
    .A3(\w[6][28] ),
    .S0(net445),
    .S1(net452),
    .X(_11406_));
 sky130_fd_sc_hd__mux4_2 _25602_ (.A0(\w[8][28] ),
    .A1(\w[12][28] ),
    .A2(\w[10][28] ),
    .A3(\w[14][28] ),
    .S0(net445),
    .S1(net452),
    .X(_11407_));
 sky130_fd_sc_hd__mux4_2 _25603_ (.A0(\w[16][28] ),
    .A1(\w[20][28] ),
    .A2(\w[18][28] ),
    .A3(\w[22][28] ),
    .S0(net445),
    .S1(net452),
    .X(_11408_));
 sky130_fd_sc_hd__mux4_2 _25604_ (.A0(\w[24][28] ),
    .A1(\w[28][28] ),
    .A2(\w[26][28] ),
    .A3(\w[30][28] ),
    .S0(net445),
    .S1(net452),
    .X(_11409_));
 sky130_fd_sc_hd__mux4_2 _25605_ (.A0(_11406_),
    .A1(_11407_),
    .A2(_11408_),
    .A3(_11409_),
    .S0(net437),
    .S1(net435),
    .X(_11410_));
 sky130_fd_sc_hd__mux4_2 _25606_ (.A0(\w[32][28] ),
    .A1(\w[36][28] ),
    .A2(\w[34][28] ),
    .A3(\w[38][28] ),
    .S0(net442),
    .S1(net450),
    .X(_11411_));
 sky130_fd_sc_hd__mux4_2 _25607_ (.A0(\w[40][28] ),
    .A1(\w[44][28] ),
    .A2(\w[42][28] ),
    .A3(\w[46][28] ),
    .S0(net442),
    .S1(net450),
    .X(_11412_));
 sky130_fd_sc_hd__mux4_2 _25608_ (.A0(\w[48][28] ),
    .A1(\w[52][28] ),
    .A2(\w[50][28] ),
    .A3(\w[54][28] ),
    .S0(net442),
    .S1(net450),
    .X(_11413_));
 sky130_fd_sc_hd__mux4_2 _25609_ (.A0(\w[56][28] ),
    .A1(\w[60][28] ),
    .A2(\w[58][28] ),
    .A3(\w[62][28] ),
    .S0(net442),
    .S1(net450),
    .X(_11414_));
 sky130_fd_sc_hd__mux4_2 _25610_ (.A0(_11411_),
    .A1(_11412_),
    .A2(_11413_),
    .A3(_11414_),
    .S0(net437),
    .S1(net435),
    .X(_11415_));
 sky130_fd_sc_hd__mux2i_4 _25611_ (.A0(_11410_),
    .A1(_11415_),
    .S(net433),
    .Y(_11416_));
 sky130_fd_sc_hd__xnor2_1 _25612_ (.A(_11346_),
    .B(_11416_),
    .Y(_11417_));
 sky130_fd_sc_hd__xnor2_1 _25613_ (.A(_11090_),
    .B(_11417_),
    .Y(_11656_));
 sky130_fd_sc_hd__mux4_2 _25614_ (.A0(\w[1][17] ),
    .A1(\w[5][17] ),
    .A2(\w[3][17] ),
    .A3(\w[7][17] ),
    .S0(net520),
    .S1(net528),
    .X(_11418_));
 sky130_fd_sc_hd__mux4_2 _25615_ (.A0(\w[9][17] ),
    .A1(\w[13][17] ),
    .A2(\w[11][17] ),
    .A3(\w[15][17] ),
    .S0(net520),
    .S1(net528),
    .X(_11419_));
 sky130_fd_sc_hd__mux4_2 _25616_ (.A0(\w[17][17] ),
    .A1(\w[21][17] ),
    .A2(\w[19][17] ),
    .A3(\w[23][17] ),
    .S0(net520),
    .S1(net528),
    .X(_11420_));
 sky130_fd_sc_hd__mux4_2 _25617_ (.A0(\w[25][17] ),
    .A1(\w[29][17] ),
    .A2(\w[27][17] ),
    .A3(\w[31][17] ),
    .S0(net520),
    .S1(net528),
    .X(_11421_));
 sky130_fd_sc_hd__mux4_2 _25618_ (.A0(_11418_),
    .A1(_11419_),
    .A2(_11420_),
    .A3(_11421_),
    .S0(net516),
    .S1(net514),
    .X(_11422_));
 sky130_fd_sc_hd__mux4_2 _25619_ (.A0(\w[33][17] ),
    .A1(\w[37][17] ),
    .A2(\w[35][17] ),
    .A3(\w[39][17] ),
    .S0(net520),
    .S1(net531),
    .X(_11423_));
 sky130_fd_sc_hd__mux4_2 _25620_ (.A0(\w[41][17] ),
    .A1(\w[45][17] ),
    .A2(\w[43][17] ),
    .A3(\w[47][17] ),
    .S0(net520),
    .S1(net531),
    .X(_11424_));
 sky130_fd_sc_hd__mux4_2 _25621_ (.A0(\w[49][17] ),
    .A1(\w[53][17] ),
    .A2(\w[51][17] ),
    .A3(\w[55][17] ),
    .S0(net520),
    .S1(net531),
    .X(_11425_));
 sky130_fd_sc_hd__mux4_2 _25622_ (.A0(\w[57][17] ),
    .A1(\w[61][17] ),
    .A2(\w[59][17] ),
    .A3(\w[63][17] ),
    .S0(net520),
    .S1(net531),
    .X(_11426_));
 sky130_fd_sc_hd__mux4_2 _25623_ (.A0(_11423_),
    .A1(_11424_),
    .A2(_11425_),
    .A3(_11426_),
    .S0(net516),
    .S1(net514),
    .X(_11427_));
 sky130_fd_sc_hd__mux2i_4 _25624_ (.A0(_11422_),
    .A1(_11427_),
    .S(net512),
    .Y(_11428_));
 sky130_fd_sc_hd__mux4_2 _25625_ (.A0(\w[1][28] ),
    .A1(\w[5][28] ),
    .A2(\w[3][28] ),
    .A3(\w[7][28] ),
    .S0(net523),
    .S1(net532),
    .X(_11429_));
 sky130_fd_sc_hd__mux4_2 _25626_ (.A0(\w[9][28] ),
    .A1(\w[13][28] ),
    .A2(\w[11][28] ),
    .A3(\w[15][28] ),
    .S0(net523),
    .S1(net532),
    .X(_11430_));
 sky130_fd_sc_hd__mux4_2 _25627_ (.A0(\w[17][28] ),
    .A1(\w[21][28] ),
    .A2(\w[19][28] ),
    .A3(\w[23][28] ),
    .S0(net523),
    .S1(net532),
    .X(_11431_));
 sky130_fd_sc_hd__mux4_2 _25628_ (.A0(\w[25][28] ),
    .A1(\w[29][28] ),
    .A2(\w[27][28] ),
    .A3(\w[31][28] ),
    .S0(net523),
    .S1(net532),
    .X(_11432_));
 sky130_fd_sc_hd__mux4_2 _25629_ (.A0(_11429_),
    .A1(_11430_),
    .A2(_11431_),
    .A3(_11432_),
    .S0(net518),
    .S1(net549),
    .X(_11433_));
 sky130_fd_sc_hd__mux4_2 _25630_ (.A0(\w[33][28] ),
    .A1(\w[37][28] ),
    .A2(\w[35][28] ),
    .A3(\w[39][28] ),
    .S0(net523),
    .S1(net528),
    .X(_11434_));
 sky130_fd_sc_hd__mux4_2 _25631_ (.A0(\w[41][28] ),
    .A1(\w[45][28] ),
    .A2(\w[43][28] ),
    .A3(\w[47][28] ),
    .S0(net523),
    .S1(net528),
    .X(_11435_));
 sky130_fd_sc_hd__mux4_2 _25632_ (.A0(\w[49][28] ),
    .A1(\w[53][28] ),
    .A2(\w[51][28] ),
    .A3(\w[55][28] ),
    .S0(net523),
    .S1(net528),
    .X(_11436_));
 sky130_fd_sc_hd__mux4_2 _25633_ (.A0(\w[57][28] ),
    .A1(\w[61][28] ),
    .A2(\w[59][28] ),
    .A3(\w[63][28] ),
    .S0(net523),
    .S1(net532),
    .X(_11437_));
 sky130_fd_sc_hd__mux4_2 _25634_ (.A0(_11434_),
    .A1(_11435_),
    .A2(_11436_),
    .A3(_11437_),
    .S0(net518),
    .S1(net549),
    .X(_11438_));
 sky130_fd_sc_hd__mux2i_4 _25635_ (.A0(_11433_),
    .A1(_11438_),
    .S(net513),
    .Y(_11439_));
 sky130_fd_sc_hd__xnor2_1 _25636_ (.A(_11428_),
    .B(_11439_),
    .Y(_11440_));
 sky130_fd_sc_hd__xnor2_1 _25637_ (.A(_11277_),
    .B(_11440_),
    .Y(_11659_));
 sky130_fd_sc_hd__mux4_2 _25638_ (.A0(\w[0][29] ),
    .A1(\w[4][29] ),
    .A2(\w[2][29] ),
    .A3(\w[6][29] ),
    .S0(net444),
    .S1(net447),
    .X(_11441_));
 sky130_fd_sc_hd__mux4_2 _25639_ (.A0(\w[8][29] ),
    .A1(\w[12][29] ),
    .A2(\w[10][29] ),
    .A3(\w[14][29] ),
    .S0(net444),
    .S1(net447),
    .X(_11442_));
 sky130_fd_sc_hd__mux4_2 _25640_ (.A0(\w[16][29] ),
    .A1(\w[20][29] ),
    .A2(\w[18][29] ),
    .A3(\w[22][29] ),
    .S0(net444),
    .S1(net447),
    .X(_11443_));
 sky130_fd_sc_hd__mux4_2 _25641_ (.A0(\w[24][29] ),
    .A1(\w[28][29] ),
    .A2(\w[26][29] ),
    .A3(\w[30][29] ),
    .S0(net444),
    .S1(net447),
    .X(_11444_));
 sky130_fd_sc_hd__mux4_2 _25642_ (.A0(_11441_),
    .A1(_11442_),
    .A2(_11443_),
    .A3(_11444_),
    .S0(net437),
    .S1(net435),
    .X(_11445_));
 sky130_fd_sc_hd__mux4_2 _25643_ (.A0(\w[32][29] ),
    .A1(\w[36][29] ),
    .A2(\w[34][29] ),
    .A3(\w[38][29] ),
    .S0(net444),
    .S1(net447),
    .X(_11446_));
 sky130_fd_sc_hd__mux4_2 _25644_ (.A0(\w[40][29] ),
    .A1(\w[44][29] ),
    .A2(\w[42][29] ),
    .A3(\w[46][29] ),
    .S0(net444),
    .S1(net447),
    .X(_11447_));
 sky130_fd_sc_hd__mux4_2 _25645_ (.A0(\w[48][29] ),
    .A1(\w[52][29] ),
    .A2(\w[50][29] ),
    .A3(\w[54][29] ),
    .S0(net444),
    .S1(net447),
    .X(_11448_));
 sky130_fd_sc_hd__mux4_2 _25646_ (.A0(\w[56][29] ),
    .A1(\w[60][29] ),
    .A2(\w[58][29] ),
    .A3(\w[62][29] ),
    .S0(net444),
    .S1(net447),
    .X(_11449_));
 sky130_fd_sc_hd__mux4_2 _25647_ (.A0(_11446_),
    .A1(_11447_),
    .A2(_11448_),
    .A3(_11449_),
    .S0(net437),
    .S1(net435),
    .X(_11450_));
 sky130_fd_sc_hd__mux2i_4 _25648_ (.A0(_11445_),
    .A1(_11450_),
    .S(\count2_1[5] ),
    .Y(_11451_));
 sky130_fd_sc_hd__xnor2_1 _25649_ (.A(_11381_),
    .B(_11451_),
    .Y(_11452_));
 sky130_fd_sc_hd__xnor2_1 _25650_ (.A(_10995_),
    .B(_11452_),
    .Y(_11664_));
 sky130_fd_sc_hd__mux4_2 _25651_ (.A0(\w[1][29] ),
    .A1(\w[5][29] ),
    .A2(\w[3][29] ),
    .A3(\w[7][29] ),
    .S0(\count15_1[2] ),
    .S1(net532),
    .X(_11453_));
 sky130_fd_sc_hd__mux4_2 _25652_ (.A0(\w[9][29] ),
    .A1(\w[13][29] ),
    .A2(\w[11][29] ),
    .A3(\w[15][29] ),
    .S0(\count15_1[2] ),
    .S1(net532),
    .X(_11454_));
 sky130_fd_sc_hd__mux4_2 _25653_ (.A0(\w[17][29] ),
    .A1(\w[21][29] ),
    .A2(\w[19][29] ),
    .A3(\w[23][29] ),
    .S0(\count15_1[2] ),
    .S1(net532),
    .X(_11455_));
 sky130_fd_sc_hd__mux4_2 _25654_ (.A0(\w[25][29] ),
    .A1(\w[29][29] ),
    .A2(\w[27][29] ),
    .A3(\w[31][29] ),
    .S0(\count15_1[2] ),
    .S1(net532),
    .X(_11456_));
 sky130_fd_sc_hd__mux4_2 _25655_ (.A0(_11453_),
    .A1(_11454_),
    .A2(_11455_),
    .A3(_11456_),
    .S0(net518),
    .S1(net549),
    .X(_11457_));
 sky130_fd_sc_hd__mux4_2 _25656_ (.A0(\w[33][29] ),
    .A1(\w[37][29] ),
    .A2(\w[35][29] ),
    .A3(\w[39][29] ),
    .S0(net522),
    .S1(\count15_1[1] ),
    .X(_11458_));
 sky130_fd_sc_hd__mux4_2 _25657_ (.A0(\w[41][29] ),
    .A1(\w[45][29] ),
    .A2(\w[43][29] ),
    .A3(\w[47][29] ),
    .S0(net522),
    .S1(\count15_1[1] ),
    .X(_11459_));
 sky130_fd_sc_hd__mux4_2 _25658_ (.A0(\w[49][29] ),
    .A1(\w[53][29] ),
    .A2(\w[51][29] ),
    .A3(\w[55][29] ),
    .S0(net523),
    .S1(\count15_1[1] ),
    .X(_11460_));
 sky130_fd_sc_hd__mux4_2 _25659_ (.A0(\w[57][29] ),
    .A1(\w[61][29] ),
    .A2(\w[59][29] ),
    .A3(\w[63][29] ),
    .S0(net523),
    .S1(\count15_1[1] ),
    .X(_11461_));
 sky130_fd_sc_hd__mux4_2 _25660_ (.A0(_11458_),
    .A1(_11459_),
    .A2(_11460_),
    .A3(_11461_),
    .S0(net518),
    .S1(net549),
    .X(_11462_));
 sky130_fd_sc_hd__mux2i_4 _25661_ (.A0(_11457_),
    .A1(_11462_),
    .S(net513),
    .Y(_11463_));
 sky130_fd_sc_hd__xnor2_1 _25662_ (.A(_11312_),
    .B(_11463_),
    .Y(_11464_));
 sky130_fd_sc_hd__xnor2_1 _25663_ (.A(_10865_),
    .B(_11464_),
    .Y(_11667_));
 sky130_fd_sc_hd__mux4_2 _25664_ (.A0(\w[0][30] ),
    .A1(\w[4][30] ),
    .A2(\w[2][30] ),
    .A3(\w[6][30] ),
    .S0(net444),
    .S1(net447),
    .X(_11465_));
 sky130_fd_sc_hd__mux4_2 _25665_ (.A0(\w[8][30] ),
    .A1(\w[12][30] ),
    .A2(\w[10][30] ),
    .A3(\w[14][30] ),
    .S0(net444),
    .S1(net447),
    .X(_11466_));
 sky130_fd_sc_hd__mux4_2 _25666_ (.A0(\w[16][30] ),
    .A1(\w[20][30] ),
    .A2(\w[18][30] ),
    .A3(\w[22][30] ),
    .S0(net444),
    .S1(net447),
    .X(_11467_));
 sky130_fd_sc_hd__mux4_2 _25667_ (.A0(\w[24][30] ),
    .A1(\w[28][30] ),
    .A2(\w[26][30] ),
    .A3(\w[30][30] ),
    .S0(net444),
    .S1(net447),
    .X(_11468_));
 sky130_fd_sc_hd__mux4_2 _25668_ (.A0(_11465_),
    .A1(_11466_),
    .A2(_11467_),
    .A3(_11468_),
    .S0(net437),
    .S1(net435),
    .X(_11469_));
 sky130_fd_sc_hd__mux4_2 _25669_ (.A0(\w[32][30] ),
    .A1(\w[36][30] ),
    .A2(\w[34][30] ),
    .A3(\w[38][30] ),
    .S0(net444),
    .S1(net447),
    .X(_11470_));
 sky130_fd_sc_hd__mux4_2 _25670_ (.A0(\w[40][30] ),
    .A1(\w[44][30] ),
    .A2(\w[42][30] ),
    .A3(\w[46][30] ),
    .S0(net444),
    .S1(net447),
    .X(_11471_));
 sky130_fd_sc_hd__mux4_2 _25671_ (.A0(\w[48][30] ),
    .A1(\w[52][30] ),
    .A2(\w[50][30] ),
    .A3(\w[54][30] ),
    .S0(net444),
    .S1(net447),
    .X(_11472_));
 sky130_fd_sc_hd__mux4_2 _25672_ (.A0(\w[56][30] ),
    .A1(\w[60][30] ),
    .A2(\w[58][30] ),
    .A3(\w[62][30] ),
    .S0(net444),
    .S1(net447),
    .X(_11473_));
 sky130_fd_sc_hd__mux4_2 _25673_ (.A0(_11470_),
    .A1(_11471_),
    .A2(_11472_),
    .A3(_11473_),
    .S0(net437),
    .S1(net435),
    .X(_11474_));
 sky130_fd_sc_hd__mux2i_4 _25674_ (.A0(_11469_),
    .A1(_11474_),
    .S(\count2_1[5] ),
    .Y(_11475_));
 sky130_fd_sc_hd__xnor2_1 _25675_ (.A(_11416_),
    .B(_11475_),
    .Y(_11476_));
 sky130_fd_sc_hd__xnor2_1 _25676_ (.A(_11071_),
    .B(_11476_),
    .Y(_11672_));
 sky130_fd_sc_hd__mux4_2 _25677_ (.A0(\w[1][30] ),
    .A1(\w[5][30] ),
    .A2(\w[3][30] ),
    .A3(\w[7][30] ),
    .S0(\count15_1[2] ),
    .S1(net532),
    .X(_11477_));
 sky130_fd_sc_hd__mux4_2 _25678_ (.A0(\w[9][30] ),
    .A1(\w[13][30] ),
    .A2(\w[11][30] ),
    .A3(\w[15][30] ),
    .S0(\count15_1[2] ),
    .S1(net532),
    .X(_11478_));
 sky130_fd_sc_hd__mux4_2 _25679_ (.A0(\w[17][30] ),
    .A1(\w[21][30] ),
    .A2(\w[19][30] ),
    .A3(\w[23][30] ),
    .S0(\count15_1[2] ),
    .S1(net532),
    .X(_11479_));
 sky130_fd_sc_hd__mux4_2 _25680_ (.A0(\w[25][30] ),
    .A1(\w[29][30] ),
    .A2(\w[27][30] ),
    .A3(\w[31][30] ),
    .S0(\count15_1[2] ),
    .S1(net532),
    .X(_11480_));
 sky130_fd_sc_hd__mux4_2 _25681_ (.A0(_11477_),
    .A1(_11478_),
    .A2(_11479_),
    .A3(_11480_),
    .S0(net518),
    .S1(net549),
    .X(_11481_));
 sky130_fd_sc_hd__mux4_2 _25682_ (.A0(\w[33][30] ),
    .A1(\w[37][30] ),
    .A2(\w[35][30] ),
    .A3(\w[39][30] ),
    .S0(net527),
    .S1(net550),
    .X(_11482_));
 sky130_fd_sc_hd__mux4_2 _25683_ (.A0(\w[41][30] ),
    .A1(\w[45][30] ),
    .A2(\w[43][30] ),
    .A3(\w[47][30] ),
    .S0(net527),
    .S1(net550),
    .X(_11483_));
 sky130_fd_sc_hd__mux4_2 _25684_ (.A0(\w[49][30] ),
    .A1(\w[53][30] ),
    .A2(\w[51][30] ),
    .A3(\w[55][30] ),
    .S0(net527),
    .S1(net550),
    .X(_11484_));
 sky130_fd_sc_hd__mux4_2 _25685_ (.A0(\w[57][30] ),
    .A1(\w[61][30] ),
    .A2(\w[59][30] ),
    .A3(\w[63][30] ),
    .S0(\count15_1[2] ),
    .S1(net550),
    .X(_11485_));
 sky130_fd_sc_hd__mux4_2 _25686_ (.A0(_11482_),
    .A1(_11483_),
    .A2(_11484_),
    .A3(_11485_),
    .S0(net518),
    .S1(net515),
    .X(_11486_));
 sky130_fd_sc_hd__mux2i_2 _25687_ (.A0(_11481_),
    .A1(_11486_),
    .S(net513),
    .Y(_11487_));
 sky130_fd_sc_hd__xnor2_1 _25688_ (.A(_11369_),
    .B(_11487_),
    .Y(_11488_));
 sky130_fd_sc_hd__xnor2_1 _25689_ (.A(_10928_),
    .B(_11488_),
    .Y(_11675_));
 sky130_fd_sc_hd__mux4_2 _25690_ (.A0(\w[0][31] ),
    .A1(\w[4][31] ),
    .A2(\w[2][31] ),
    .A3(\w[6][31] ),
    .S0(net442),
    .S1(net450),
    .X(_11489_));
 sky130_fd_sc_hd__mux4_2 _25691_ (.A0(\w[8][31] ),
    .A1(\w[12][31] ),
    .A2(\w[10][31] ),
    .A3(\w[14][31] ),
    .S0(net442),
    .S1(net450),
    .X(_11490_));
 sky130_fd_sc_hd__mux4_2 _25692_ (.A0(\w[16][31] ),
    .A1(\w[20][31] ),
    .A2(\w[18][31] ),
    .A3(\w[22][31] ),
    .S0(net441),
    .S1(net449),
    .X(_11491_));
 sky130_fd_sc_hd__mux4_2 _25693_ (.A0(\w[24][31] ),
    .A1(\w[28][31] ),
    .A2(\w[26][31] ),
    .A3(\w[30][31] ),
    .S0(net441),
    .S1(net449),
    .X(_11492_));
 sky130_fd_sc_hd__mux4_2 _25694_ (.A0(_11489_),
    .A1(_11490_),
    .A2(_11491_),
    .A3(_11492_),
    .S0(net438),
    .S1(net434),
    .X(_11493_));
 sky130_fd_sc_hd__mux4_2 _25695_ (.A0(\w[32][31] ),
    .A1(\w[36][31] ),
    .A2(\w[34][31] ),
    .A3(\w[38][31] ),
    .S0(net441),
    .S1(net449),
    .X(_11494_));
 sky130_fd_sc_hd__mux4_2 _25696_ (.A0(\w[40][31] ),
    .A1(\w[44][31] ),
    .A2(\w[42][31] ),
    .A3(\w[46][31] ),
    .S0(net441),
    .S1(net449),
    .X(_11495_));
 sky130_fd_sc_hd__mux4_2 _25697_ (.A0(\w[48][31] ),
    .A1(\w[52][31] ),
    .A2(\w[50][31] ),
    .A3(\w[54][31] ),
    .S0(net441),
    .S1(net449),
    .X(_11496_));
 sky130_fd_sc_hd__mux4_2 _25698_ (.A0(\w[56][31] ),
    .A1(\w[60][31] ),
    .A2(\w[58][31] ),
    .A3(\w[62][31] ),
    .S0(net443),
    .S1(net451),
    .X(_11497_));
 sky130_fd_sc_hd__mux4_2 _25699_ (.A0(_11494_),
    .A1(_11495_),
    .A2(_11496_),
    .A3(_11497_),
    .S0(net438),
    .S1(net434),
    .X(_11498_));
 sky130_fd_sc_hd__mux2i_4 _25700_ (.A0(_11493_),
    .A1(_11498_),
    .S(net432),
    .Y(_11499_));
 sky130_fd_sc_hd__xnor2_1 _25701_ (.A(_11451_),
    .B(_11499_),
    .Y(_11500_));
 sky130_fd_sc_hd__xnor2_1 _25702_ (.A(_11158_),
    .B(_11500_),
    .Y(_11680_));
 sky130_fd_sc_hd__mux4_2 _25703_ (.A0(\w[1][31] ),
    .A1(\w[5][31] ),
    .A2(\w[3][31] ),
    .A3(\w[7][31] ),
    .S0(net520),
    .S1(net528),
    .X(_11501_));
 sky130_fd_sc_hd__mux4_2 _25704_ (.A0(\w[9][31] ),
    .A1(\w[13][31] ),
    .A2(\w[11][31] ),
    .A3(\w[15][31] ),
    .S0(net520),
    .S1(net528),
    .X(_11502_));
 sky130_fd_sc_hd__mux4_2 _25705_ (.A0(\w[17][31] ),
    .A1(\w[21][31] ),
    .A2(\w[19][31] ),
    .A3(\w[23][31] ),
    .S0(net520),
    .S1(net528),
    .X(_11503_));
 sky130_fd_sc_hd__mux4_2 _25706_ (.A0(\w[25][31] ),
    .A1(\w[29][31] ),
    .A2(\w[27][31] ),
    .A3(\w[31][31] ),
    .S0(net520),
    .S1(net528),
    .X(_11504_));
 sky130_fd_sc_hd__mux4_2 _25707_ (.A0(_11501_),
    .A1(_11502_),
    .A2(_11503_),
    .A3(_11504_),
    .S0(net516),
    .S1(net514),
    .X(_11505_));
 sky130_fd_sc_hd__mux4_2 _25708_ (.A0(\w[33][31] ),
    .A1(\w[37][31] ),
    .A2(\w[35][31] ),
    .A3(\w[39][31] ),
    .S0(net519),
    .S1(net528),
    .X(_11506_));
 sky130_fd_sc_hd__mux4_2 _25709_ (.A0(\w[41][31] ),
    .A1(\w[45][31] ),
    .A2(\w[43][31] ),
    .A3(\w[47][31] ),
    .S0(net519),
    .S1(net528),
    .X(_11507_));
 sky130_fd_sc_hd__mux4_2 _25710_ (.A0(\w[49][31] ),
    .A1(\w[53][31] ),
    .A2(\w[51][31] ),
    .A3(\w[55][31] ),
    .S0(net519),
    .S1(net528),
    .X(_11508_));
 sky130_fd_sc_hd__mux4_2 _25711_ (.A0(\w[57][31] ),
    .A1(\w[61][31] ),
    .A2(\w[59][31] ),
    .A3(\w[63][31] ),
    .S0(net519),
    .S1(net528),
    .X(_11509_));
 sky130_fd_sc_hd__mux4_2 _25712_ (.A0(_11506_),
    .A1(_11507_),
    .A2(_11508_),
    .A3(_11509_),
    .S0(net518),
    .S1(net549),
    .X(_11510_));
 sky130_fd_sc_hd__mux2i_4 _25713_ (.A0(_11505_),
    .A1(_11510_),
    .S(net512),
    .Y(_11511_));
 sky130_fd_sc_hd__xnor2_1 _25714_ (.A(_11404_),
    .B(_11511_),
    .Y(_11512_));
 sky130_fd_sc_hd__xnor2_1 _25715_ (.A(_11022_),
    .B(_11512_),
    .Y(_11683_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_286 ();
 sky130_fd_sc_hd__mux4_2 _25718_ (.A0(\w[0][0] ),
    .A1(\w[4][0] ),
    .A2(\w[2][0] ),
    .A3(\w[6][0] ),
    .S0(net439),
    .S1(net448),
    .X(_11515_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_284 ();
 sky130_fd_sc_hd__mux4_2 _25721_ (.A0(\w[8][0] ),
    .A1(\w[12][0] ),
    .A2(\w[10][0] ),
    .A3(\w[14][0] ),
    .S0(net439),
    .S1(net448),
    .X(_11518_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_282 ();
 sky130_fd_sc_hd__mux4_2 _25724_ (.A0(\w[16][0] ),
    .A1(\w[20][0] ),
    .A2(\w[18][0] ),
    .A3(\w[22][0] ),
    .S0(net439),
    .S1(net448),
    .X(_11521_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_280 ();
 sky130_fd_sc_hd__mux4_2 _25727_ (.A0(\w[24][0] ),
    .A1(\w[28][0] ),
    .A2(\w[26][0] ),
    .A3(\w[30][0] ),
    .S0(net439),
    .S1(net448),
    .X(_11524_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_278 ();
 sky130_fd_sc_hd__mux4_2 _25730_ (.A0(_11515_),
    .A1(_11518_),
    .A2(_11521_),
    .A3(_11524_),
    .S0(net436),
    .S1(net434),
    .X(_11527_));
 sky130_fd_sc_hd__mux4_2 _25731_ (.A0(\w[32][0] ),
    .A1(\w[36][0] ),
    .A2(\w[34][0] ),
    .A3(\w[38][0] ),
    .S0(net441),
    .S1(net449),
    .X(_11528_));
 sky130_fd_sc_hd__mux4_2 _25732_ (.A0(\w[40][0] ),
    .A1(\w[44][0] ),
    .A2(\w[42][0] ),
    .A3(\w[46][0] ),
    .S0(net441),
    .S1(net449),
    .X(_11529_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_276 ();
 sky130_fd_sc_hd__mux4_2 _25735_ (.A0(\w[48][0] ),
    .A1(\w[52][0] ),
    .A2(\w[50][0] ),
    .A3(\w[54][0] ),
    .S0(net441),
    .S1(net449),
    .X(_11532_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_274 ();
 sky130_fd_sc_hd__mux4_2 _25738_ (.A0(\w[56][0] ),
    .A1(\w[60][0] ),
    .A2(\w[58][0] ),
    .A3(\w[62][0] ),
    .S0(net441),
    .S1(net449),
    .X(_11535_));
 sky130_fd_sc_hd__mux4_2 _25739_ (.A0(_11528_),
    .A1(_11529_),
    .A2(_11532_),
    .A3(_11535_),
    .S0(net436),
    .S1(net434),
    .X(_11536_));
 sky130_fd_sc_hd__mux2i_4 _25740_ (.A0(_11527_),
    .A1(_11536_),
    .S(net432),
    .Y(_11537_));
 sky130_fd_sc_hd__xnor2_1 _25741_ (.A(_11475_),
    .B(_11537_),
    .Y(_11538_));
 sky130_fd_sc_hd__xnor2_1 _25742_ (.A(_11207_),
    .B(_11538_),
    .Y(_11688_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_272 ();
 sky130_fd_sc_hd__mux4_2 _25745_ (.A0(\w[1][0] ),
    .A1(\w[5][0] ),
    .A2(\w[3][0] ),
    .A3(\w[7][0] ),
    .S0(net521),
    .S1(net528),
    .X(_11541_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_270 ();
 sky130_fd_sc_hd__mux4_2 _25748_ (.A0(\w[9][0] ),
    .A1(\w[13][0] ),
    .A2(\w[11][0] ),
    .A3(\w[15][0] ),
    .S0(net521),
    .S1(net528),
    .X(_11544_));
 sky130_fd_sc_hd__mux4_2 _25749_ (.A0(\w[17][0] ),
    .A1(\w[21][0] ),
    .A2(\w[19][0] ),
    .A3(\w[23][0] ),
    .S0(net521),
    .S1(net528),
    .X(_11545_));
 sky130_fd_sc_hd__mux4_2 _25750_ (.A0(\w[25][0] ),
    .A1(\w[29][0] ),
    .A2(\w[27][0] ),
    .A3(\w[31][0] ),
    .S0(net521),
    .S1(net528),
    .X(_11546_));
 sky130_fd_sc_hd__mux4_2 _25751_ (.A0(_11541_),
    .A1(_11544_),
    .A2(_11545_),
    .A3(_11546_),
    .S0(net516),
    .S1(net514),
    .X(_11547_));
 sky130_fd_sc_hd__mux4_2 _25752_ (.A0(\w[33][0] ),
    .A1(\w[37][0] ),
    .A2(\w[35][0] ),
    .A3(\w[39][0] ),
    .S0(net521),
    .S1(net531),
    .X(_11548_));
 sky130_fd_sc_hd__mux4_2 _25753_ (.A0(\w[41][0] ),
    .A1(\w[45][0] ),
    .A2(\w[43][0] ),
    .A3(\w[47][0] ),
    .S0(net521),
    .S1(net531),
    .X(_11549_));
 sky130_fd_sc_hd__mux4_2 _25754_ (.A0(\w[49][0] ),
    .A1(\w[53][0] ),
    .A2(\w[51][0] ),
    .A3(\w[55][0] ),
    .S0(net521),
    .S1(net531),
    .X(_11550_));
 sky130_fd_sc_hd__mux4_2 _25755_ (.A0(\w[57][0] ),
    .A1(\w[61][0] ),
    .A2(\w[59][0] ),
    .A3(\w[63][0] ),
    .S0(net521),
    .S1(net531),
    .X(_11551_));
 sky130_fd_sc_hd__mux4_2 _25756_ (.A0(_11548_),
    .A1(_11549_),
    .A2(_11550_),
    .A3(_11551_),
    .S0(net516),
    .S1(net514),
    .X(_11552_));
 sky130_fd_sc_hd__mux2i_4 _25757_ (.A0(_11547_),
    .A1(_11552_),
    .S(net512),
    .Y(_11553_));
 sky130_fd_sc_hd__xnor2_1 _25758_ (.A(_11428_),
    .B(_11553_),
    .Y(_11554_));
 sky130_fd_sc_hd__xnor2_1 _25759_ (.A(_11117_),
    .B(_11554_),
    .Y(_11691_));
 sky130_fd_sc_hd__mux4_2 _25760_ (.A0(\w[0][1] ),
    .A1(\w[4][1] ),
    .A2(\w[2][1] ),
    .A3(\w[6][1] ),
    .S0(net439),
    .S1(net448),
    .X(_11555_));
 sky130_fd_sc_hd__mux4_2 _25761_ (.A0(\w[8][1] ),
    .A1(\w[12][1] ),
    .A2(\w[10][1] ),
    .A3(\w[14][1] ),
    .S0(net439),
    .S1(net448),
    .X(_11556_));
 sky130_fd_sc_hd__mux4_2 _25762_ (.A0(\w[16][1] ),
    .A1(\w[20][1] ),
    .A2(\w[18][1] ),
    .A3(\w[22][1] ),
    .S0(net439),
    .S1(net448),
    .X(_11557_));
 sky130_fd_sc_hd__mux4_2 _25763_ (.A0(\w[24][1] ),
    .A1(\w[28][1] ),
    .A2(\w[26][1] ),
    .A3(\w[30][1] ),
    .S0(net439),
    .S1(net448),
    .X(_11558_));
 sky130_fd_sc_hd__mux4_2 _25764_ (.A0(_11555_),
    .A1(_11556_),
    .A2(_11557_),
    .A3(_11558_),
    .S0(net436),
    .S1(net434),
    .X(_11559_));
 sky130_fd_sc_hd__mux4_2 _25765_ (.A0(\w[32][1] ),
    .A1(\w[36][1] ),
    .A2(\w[34][1] ),
    .A3(\w[38][1] ),
    .S0(net443),
    .S1(net451),
    .X(_11560_));
 sky130_fd_sc_hd__mux4_2 _25766_ (.A0(\w[40][1] ),
    .A1(\w[44][1] ),
    .A2(\w[42][1] ),
    .A3(\w[46][1] ),
    .S0(net443),
    .S1(net451),
    .X(_11561_));
 sky130_fd_sc_hd__mux4_2 _25767_ (.A0(\w[48][1] ),
    .A1(\w[52][1] ),
    .A2(\w[50][1] ),
    .A3(\w[54][1] ),
    .S0(net443),
    .S1(net451),
    .X(_11562_));
 sky130_fd_sc_hd__mux4_2 _25768_ (.A0(\w[56][1] ),
    .A1(\w[60][1] ),
    .A2(\w[58][1] ),
    .A3(\w[62][1] ),
    .S0(net443),
    .S1(net451),
    .X(_11563_));
 sky130_fd_sc_hd__mux4_2 _25769_ (.A0(_11560_),
    .A1(_11561_),
    .A2(_11562_),
    .A3(_11563_),
    .S0(net436),
    .S1(net434),
    .X(_11564_));
 sky130_fd_sc_hd__mux2i_4 _25770_ (.A0(_11559_),
    .A1(_11564_),
    .S(net432),
    .Y(_11565_));
 sky130_fd_sc_hd__xnor2_1 _25771_ (.A(_11499_),
    .B(_11565_),
    .Y(_11566_));
 sky130_fd_sc_hd__xnor2_1 _25772_ (.A(_11254_),
    .B(_11566_),
    .Y(_11696_));
 sky130_fd_sc_hd__mux4_2 _25773_ (.A0(\w[1][1] ),
    .A1(\w[5][1] ),
    .A2(\w[3][1] ),
    .A3(\w[7][1] ),
    .S0(net520),
    .S1(net528),
    .X(_11567_));
 sky130_fd_sc_hd__mux4_2 _25774_ (.A0(\w[9][1] ),
    .A1(\w[13][1] ),
    .A2(\w[11][1] ),
    .A3(\w[15][1] ),
    .S0(net520),
    .S1(net528),
    .X(_11568_));
 sky130_fd_sc_hd__mux4_2 _25775_ (.A0(\w[17][1] ),
    .A1(\w[21][1] ),
    .A2(\w[19][1] ),
    .A3(\w[23][1] ),
    .S0(net520),
    .S1(net528),
    .X(_11569_));
 sky130_fd_sc_hd__mux4_2 _25776_ (.A0(\w[25][1] ),
    .A1(\w[29][1] ),
    .A2(\w[27][1] ),
    .A3(\w[31][1] ),
    .S0(net520),
    .S1(net528),
    .X(_11570_));
 sky130_fd_sc_hd__mux4_2 _25777_ (.A0(_11567_),
    .A1(_11568_),
    .A2(_11569_),
    .A3(_11570_),
    .S0(net516),
    .S1(net514),
    .X(_11571_));
 sky130_fd_sc_hd__mux4_2 _25778_ (.A0(\w[33][1] ),
    .A1(\w[37][1] ),
    .A2(\w[35][1] ),
    .A3(\w[39][1] ),
    .S0(net519),
    .S1(net528),
    .X(_11572_));
 sky130_fd_sc_hd__mux4_2 _25779_ (.A0(\w[41][1] ),
    .A1(\w[45][1] ),
    .A2(\w[43][1] ),
    .A3(\w[47][1] ),
    .S0(net519),
    .S1(net528),
    .X(_11573_));
 sky130_fd_sc_hd__mux4_2 _25780_ (.A0(\w[49][1] ),
    .A1(\w[53][1] ),
    .A2(\w[51][1] ),
    .A3(\w[55][1] ),
    .S0(net519),
    .S1(net528),
    .X(_11574_));
 sky130_fd_sc_hd__mux4_2 _25781_ (.A0(\w[57][1] ),
    .A1(\w[61][1] ),
    .A2(\w[59][1] ),
    .A3(\w[63][1] ),
    .S0(net519),
    .S1(net528),
    .X(_02570_));
 sky130_fd_sc_hd__mux4_2 _25782_ (.A0(_11572_),
    .A1(_11573_),
    .A2(_11574_),
    .A3(_02570_),
    .S0(net516),
    .S1(net514),
    .X(_02571_));
 sky130_fd_sc_hd__mux2i_4 _25783_ (.A0(_11571_),
    .A1(_02571_),
    .S(net512),
    .Y(_02572_));
 sky130_fd_sc_hd__xnor2_1 _25784_ (.A(_11172_),
    .B(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__xnor2_1 _25785_ (.A(_10865_),
    .B(_02573_),
    .Y(_11699_));
 sky130_fd_sc_hd__mux4_2 _25786_ (.A0(\w[0][2] ),
    .A1(\w[4][2] ),
    .A2(\w[2][2] ),
    .A3(\w[6][2] ),
    .S0(net444),
    .S1(net447),
    .X(_02574_));
 sky130_fd_sc_hd__mux4_2 _25787_ (.A0(\w[8][2] ),
    .A1(\w[12][2] ),
    .A2(\w[10][2] ),
    .A3(\w[14][2] ),
    .S0(net444),
    .S1(net447),
    .X(_02575_));
 sky130_fd_sc_hd__mux4_2 _25788_ (.A0(\w[16][2] ),
    .A1(\w[20][2] ),
    .A2(\w[18][2] ),
    .A3(\w[22][2] ),
    .S0(net444),
    .S1(net447),
    .X(_02576_));
 sky130_fd_sc_hd__mux4_2 _25789_ (.A0(\w[24][2] ),
    .A1(\w[28][2] ),
    .A2(\w[26][2] ),
    .A3(\w[30][2] ),
    .S0(net444),
    .S1(net447),
    .X(_02577_));
 sky130_fd_sc_hd__mux4_2 _25790_ (.A0(_02574_),
    .A1(_02575_),
    .A2(_02576_),
    .A3(_02577_),
    .S0(net437),
    .S1(net435),
    .X(_02578_));
 sky130_fd_sc_hd__mux4_2 _25791_ (.A0(\w[32][2] ),
    .A1(\w[36][2] ),
    .A2(\w[34][2] ),
    .A3(\w[38][2] ),
    .S0(net445),
    .S1(net452),
    .X(_02579_));
 sky130_fd_sc_hd__mux4_2 _25792_ (.A0(\w[40][2] ),
    .A1(\w[44][2] ),
    .A2(\w[42][2] ),
    .A3(\w[46][2] ),
    .S0(net445),
    .S1(net452),
    .X(_02580_));
 sky130_fd_sc_hd__mux4_2 _25793_ (.A0(\w[48][2] ),
    .A1(\w[52][2] ),
    .A2(\w[50][2] ),
    .A3(\w[54][2] ),
    .S0(net445),
    .S1(net452),
    .X(_02581_));
 sky130_fd_sc_hd__mux4_2 _25794_ (.A0(\w[56][2] ),
    .A1(\w[60][2] ),
    .A2(\w[58][2] ),
    .A3(\w[62][2] ),
    .S0(net445),
    .S1(net452),
    .X(_02582_));
 sky130_fd_sc_hd__mux4_2 _25795_ (.A0(_02579_),
    .A1(_02580_),
    .A2(_02581_),
    .A3(_02582_),
    .S0(net437),
    .S1(net435),
    .X(_02583_));
 sky130_fd_sc_hd__mux2i_4 _25796_ (.A0(_02578_),
    .A1(_02583_),
    .S(net433),
    .Y(_02584_));
 sky130_fd_sc_hd__xnor2_1 _25797_ (.A(_11537_),
    .B(_02584_),
    .Y(_02585_));
 sky130_fd_sc_hd__xnor2_1 _25798_ (.A(_11289_),
    .B(_02585_),
    .Y(_11704_));
 sky130_fd_sc_hd__mux4_2 _25799_ (.A0(\w[1][2] ),
    .A1(\w[5][2] ),
    .A2(\w[3][2] ),
    .A3(\w[7][2] ),
    .S0(net521),
    .S1(net531),
    .X(_02586_));
 sky130_fd_sc_hd__mux4_2 _25800_ (.A0(\w[9][2] ),
    .A1(\w[13][2] ),
    .A2(\w[11][2] ),
    .A3(\w[15][2] ),
    .S0(net521),
    .S1(net531),
    .X(_02587_));
 sky130_fd_sc_hd__mux4_2 _25801_ (.A0(\w[17][2] ),
    .A1(\w[21][2] ),
    .A2(\w[19][2] ),
    .A3(\w[23][2] ),
    .S0(net521),
    .S1(net531),
    .X(_02588_));
 sky130_fd_sc_hd__mux4_2 _25802_ (.A0(\w[25][2] ),
    .A1(\w[29][2] ),
    .A2(\w[27][2] ),
    .A3(\w[31][2] ),
    .S0(net521),
    .S1(net531),
    .X(_02589_));
 sky130_fd_sc_hd__mux4_2 _25803_ (.A0(_02586_),
    .A1(_02587_),
    .A2(_02588_),
    .A3(_02589_),
    .S0(net516),
    .S1(net514),
    .X(_02590_));
 sky130_fd_sc_hd__mux4_2 _25804_ (.A0(\w[33][2] ),
    .A1(\w[37][2] ),
    .A2(\w[35][2] ),
    .A3(\w[39][2] ),
    .S0(net522),
    .S1(net531),
    .X(_02591_));
 sky130_fd_sc_hd__mux4_2 _25805_ (.A0(\w[41][2] ),
    .A1(\w[45][2] ),
    .A2(\w[43][2] ),
    .A3(\w[47][2] ),
    .S0(net522),
    .S1(net531),
    .X(_02592_));
 sky130_fd_sc_hd__mux4_2 _25806_ (.A0(\w[49][2] ),
    .A1(\w[53][2] ),
    .A2(\w[51][2] ),
    .A3(\w[55][2] ),
    .S0(net522),
    .S1(net531),
    .X(_02593_));
 sky130_fd_sc_hd__mux4_2 _25807_ (.A0(\w[57][2] ),
    .A1(\w[61][2] ),
    .A2(\w[59][2] ),
    .A3(\w[63][2] ),
    .S0(net522),
    .S1(net529),
    .X(_02594_));
 sky130_fd_sc_hd__mux4_2 _25808_ (.A0(_02591_),
    .A1(_02592_),
    .A2(_02593_),
    .A3(_02594_),
    .S0(net516),
    .S1(net514),
    .X(_02595_));
 sky130_fd_sc_hd__mux2i_4 _25809_ (.A0(_02590_),
    .A1(_02595_),
    .S(net512),
    .Y(_02596_));
 sky130_fd_sc_hd__xnor2_1 _25810_ (.A(_11220_),
    .B(_02596_),
    .Y(_02597_));
 sky130_fd_sc_hd__xnor2_1 _25811_ (.A(_10928_),
    .B(_02597_),
    .Y(_11707_));
 sky130_fd_sc_hd__mux4_2 _25812_ (.A0(\w[0][3] ),
    .A1(\w[4][3] ),
    .A2(\w[2][3] ),
    .A3(\w[6][3] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_02598_));
 sky130_fd_sc_hd__mux4_2 _25813_ (.A0(\w[8][3] ),
    .A1(\w[12][3] ),
    .A2(\w[10][3] ),
    .A3(\w[14][3] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_02599_));
 sky130_fd_sc_hd__mux4_2 _25814_ (.A0(\w[16][3] ),
    .A1(\w[20][3] ),
    .A2(\w[18][3] ),
    .A3(\w[22][3] ),
    .S0(\count2_1[2] ),
    .S1(\count2_1[1] ),
    .X(_02600_));
 sky130_fd_sc_hd__mux4_2 _25815_ (.A0(\w[24][3] ),
    .A1(\w[28][3] ),
    .A2(\w[26][3] ),
    .A3(\w[30][3] ),
    .S0(\count2_1[2] ),
    .S1(net1093),
    .X(_02601_));
 sky130_fd_sc_hd__mux4_2 _25816_ (.A0(_02598_),
    .A1(_02599_),
    .A2(_02600_),
    .A3(_02601_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_02602_));
 sky130_fd_sc_hd__mux4_2 _25817_ (.A0(\w[32][3] ),
    .A1(\w[36][3] ),
    .A2(\w[34][3] ),
    .A3(\w[38][3] ),
    .S0(\count2_1[2] ),
    .S1(net1093),
    .X(_02603_));
 sky130_fd_sc_hd__mux4_2 _25818_ (.A0(\w[40][3] ),
    .A1(\w[44][3] ),
    .A2(\w[42][3] ),
    .A3(\w[46][3] ),
    .S0(\count2_1[2] ),
    .S1(net1093),
    .X(_02604_));
 sky130_fd_sc_hd__mux4_2 _25819_ (.A0(\w[48][3] ),
    .A1(\w[52][3] ),
    .A2(\w[50][3] ),
    .A3(\w[54][3] ),
    .S0(\count2_1[2] ),
    .S1(net1093),
    .X(_02605_));
 sky130_fd_sc_hd__mux4_2 _25820_ (.A0(\w[56][3] ),
    .A1(\w[60][3] ),
    .A2(\w[58][3] ),
    .A3(\w[62][3] ),
    .S0(\count2_1[2] ),
    .S1(net452),
    .X(_02606_));
 sky130_fd_sc_hd__mux4_2 _25821_ (.A0(_02603_),
    .A1(_02604_),
    .A2(_02605_),
    .A3(_02606_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_02607_));
 sky130_fd_sc_hd__mux2i_4 _25822_ (.A0(_02602_),
    .A1(_02607_),
    .S(\count2_1[5] ),
    .Y(_02608_));
 sky130_fd_sc_hd__xnor2_1 _25823_ (.A(_11565_),
    .B(_02608_),
    .Y(_02609_));
 sky130_fd_sc_hd__xnor2_1 _25824_ (.A(_11346_),
    .B(_02609_),
    .Y(_11712_));
 sky130_fd_sc_hd__xnor2_1 _25825_ (.A(_11022_),
    .B(_11266_),
    .Y(_02610_));
 sky130_fd_sc_hd__xnor2_1 _25826_ (.A(_10833_),
    .B(_02610_),
    .Y(_11715_));
 sky130_fd_sc_hd__mux4_2 _25827_ (.A0(\w[0][4] ),
    .A1(\w[4][4] ),
    .A2(\w[2][4] ),
    .A3(\w[6][4] ),
    .S0(net444),
    .S1(net447),
    .X(_02611_));
 sky130_fd_sc_hd__mux4_2 _25828_ (.A0(\w[8][4] ),
    .A1(\w[12][4] ),
    .A2(\w[10][4] ),
    .A3(\w[14][4] ),
    .S0(net444),
    .S1(net447),
    .X(_02612_));
 sky130_fd_sc_hd__mux4_2 _25829_ (.A0(\w[16][4] ),
    .A1(\w[20][4] ),
    .A2(\w[18][4] ),
    .A3(\w[22][4] ),
    .S0(net444),
    .S1(net447),
    .X(_02613_));
 sky130_fd_sc_hd__mux4_2 _25830_ (.A0(\w[24][4] ),
    .A1(\w[28][4] ),
    .A2(\w[26][4] ),
    .A3(\w[30][4] ),
    .S0(net444),
    .S1(net447),
    .X(_02614_));
 sky130_fd_sc_hd__mux4_2 _25831_ (.A0(_02611_),
    .A1(_02612_),
    .A2(_02613_),
    .A3(_02614_),
    .S0(net437),
    .S1(net435),
    .X(_02615_));
 sky130_fd_sc_hd__mux4_2 _25832_ (.A0(\w[32][4] ),
    .A1(\w[36][4] ),
    .A2(\w[34][4] ),
    .A3(\w[38][4] ),
    .S0(net444),
    .S1(net447),
    .X(_02616_));
 sky130_fd_sc_hd__mux4_2 _25833_ (.A0(\w[40][4] ),
    .A1(\w[44][4] ),
    .A2(\w[42][4] ),
    .A3(\w[46][4] ),
    .S0(net446),
    .S1(net447),
    .X(_02617_));
 sky130_fd_sc_hd__mux4_2 _25834_ (.A0(\w[48][4] ),
    .A1(\w[52][4] ),
    .A2(\w[50][4] ),
    .A3(\w[54][4] ),
    .S0(net446),
    .S1(net447),
    .X(_02618_));
 sky130_fd_sc_hd__mux4_2 _25835_ (.A0(\w[56][4] ),
    .A1(\w[60][4] ),
    .A2(\w[58][4] ),
    .A3(\w[62][4] ),
    .S0(net446),
    .S1(net447),
    .X(_02619_));
 sky130_fd_sc_hd__mux4_2 _25836_ (.A0(_02616_),
    .A1(_02617_),
    .A2(_02618_),
    .A3(_02619_),
    .S0(net437),
    .S1(net435),
    .X(_02620_));
 sky130_fd_sc_hd__mux2i_4 _25837_ (.A0(_02615_),
    .A1(_02620_),
    .S(\count2_1[5] ),
    .Y(_02621_));
 sky130_fd_sc_hd__xnor2_1 _25838_ (.A(_02584_),
    .B(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__xnor2_1 _25839_ (.A(_11381_),
    .B(_02622_),
    .Y(_11720_));
 sky130_fd_sc_hd__xnor2_1 _25840_ (.A(_11117_),
    .B(_11323_),
    .Y(_02623_));
 sky130_fd_sc_hd__xnor2_1 _25841_ (.A(_10905_),
    .B(_02623_),
    .Y(_11723_));
 sky130_fd_sc_hd__mux4_2 _25842_ (.A0(\w[0][5] ),
    .A1(\w[4][5] ),
    .A2(\w[2][5] ),
    .A3(\w[6][5] ),
    .S0(net446),
    .S1(net447),
    .X(_02624_));
 sky130_fd_sc_hd__mux4_2 _25843_ (.A0(\w[8][5] ),
    .A1(\w[12][5] ),
    .A2(\w[10][5] ),
    .A3(\w[14][5] ),
    .S0(net446),
    .S1(net447),
    .X(_02625_));
 sky130_fd_sc_hd__mux4_2 _25844_ (.A0(\w[16][5] ),
    .A1(\w[20][5] ),
    .A2(\w[18][5] ),
    .A3(\w[22][5] ),
    .S0(net446),
    .S1(net447),
    .X(_02626_));
 sky130_fd_sc_hd__mux4_2 _25845_ (.A0(\w[24][5] ),
    .A1(\w[28][5] ),
    .A2(\w[26][5] ),
    .A3(\w[30][5] ),
    .S0(net446),
    .S1(net447),
    .X(_02627_));
 sky130_fd_sc_hd__mux4_2 _25846_ (.A0(_02624_),
    .A1(_02625_),
    .A2(_02626_),
    .A3(_02627_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_02628_));
 sky130_fd_sc_hd__mux4_2 _25847_ (.A0(\w[32][5] ),
    .A1(\w[36][5] ),
    .A2(\w[34][5] ),
    .A3(\w[38][5] ),
    .S0(net446),
    .S1(net447),
    .X(_02629_));
 sky130_fd_sc_hd__mux4_2 _25848_ (.A0(\w[40][5] ),
    .A1(\w[44][5] ),
    .A2(\w[42][5] ),
    .A3(\w[46][5] ),
    .S0(net446),
    .S1(net447),
    .X(_02630_));
 sky130_fd_sc_hd__mux4_2 _25849_ (.A0(\w[48][5] ),
    .A1(\w[52][5] ),
    .A2(\w[50][5] ),
    .A3(\w[54][5] ),
    .S0(net446),
    .S1(net447),
    .X(_02631_));
 sky130_fd_sc_hd__mux4_2 _25850_ (.A0(\w[56][5] ),
    .A1(\w[60][5] ),
    .A2(\w[58][5] ),
    .A3(\w[62][5] ),
    .S0(net446),
    .S1(net447),
    .X(_02632_));
 sky130_fd_sc_hd__mux4_2 _25851_ (.A0(_02629_),
    .A1(_02630_),
    .A2(_02631_),
    .A3(_02632_),
    .S0(net437),
    .S1(net435),
    .X(_02633_));
 sky130_fd_sc_hd__mux2i_4 _25852_ (.A0(_02628_),
    .A1(_02633_),
    .S(\count2_1[5] ),
    .Y(_02634_));
 sky130_fd_sc_hd__xnor2_1 _25853_ (.A(_02608_),
    .B(_02634_),
    .Y(_02635_));
 sky130_fd_sc_hd__xnor2_1 _25854_ (.A(_11416_),
    .B(_02635_),
    .Y(_11728_));
 sky130_fd_sc_hd__xnor2_1 _25855_ (.A(_11172_),
    .B(_11358_),
    .Y(_02636_));
 sky130_fd_sc_hd__xnor2_2 _25856_ (.A(_11034_),
    .B(_02636_),
    .Y(_11731_));
 sky130_fd_sc_hd__mux4_2 _25857_ (.A0(\w[0][6] ),
    .A1(\w[4][6] ),
    .A2(\w[2][6] ),
    .A3(\w[6][6] ),
    .S0(net446),
    .S1(net447),
    .X(_02637_));
 sky130_fd_sc_hd__mux4_2 _25858_ (.A0(\w[8][6] ),
    .A1(\w[12][6] ),
    .A2(\w[10][6] ),
    .A3(\w[14][6] ),
    .S0(net446),
    .S1(net447),
    .X(_02638_));
 sky130_fd_sc_hd__mux4_2 _25859_ (.A0(\w[16][6] ),
    .A1(\w[20][6] ),
    .A2(\w[18][6] ),
    .A3(\w[22][6] ),
    .S0(net446),
    .S1(net447),
    .X(_02639_));
 sky130_fd_sc_hd__mux4_2 _25860_ (.A0(\w[24][6] ),
    .A1(\w[28][6] ),
    .A2(\w[26][6] ),
    .A3(\w[30][6] ),
    .S0(net446),
    .S1(net447),
    .X(_02640_));
 sky130_fd_sc_hd__mux4_2 _25861_ (.A0(_02637_),
    .A1(_02638_),
    .A2(_02639_),
    .A3(_02640_),
    .S0(\count2_1[3] ),
    .S1(\count2_1[4] ),
    .X(_02641_));
 sky130_fd_sc_hd__mux4_2 _25862_ (.A0(\w[32][6] ),
    .A1(\w[36][6] ),
    .A2(\w[34][6] ),
    .A3(\w[38][6] ),
    .S0(net446),
    .S1(net1093),
    .X(_02642_));
 sky130_fd_sc_hd__mux4_2 _25863_ (.A0(\w[40][6] ),
    .A1(\w[44][6] ),
    .A2(\w[42][6] ),
    .A3(\w[46][6] ),
    .S0(net446),
    .S1(net1093),
    .X(_02643_));
 sky130_fd_sc_hd__mux4_2 _25864_ (.A0(\w[48][6] ),
    .A1(\w[52][6] ),
    .A2(\w[50][6] ),
    .A3(\w[54][6] ),
    .S0(net446),
    .S1(net1093),
    .X(_02644_));
 sky130_fd_sc_hd__mux4_2 _25865_ (.A0(\w[56][6] ),
    .A1(\w[60][6] ),
    .A2(\w[58][6] ),
    .A3(\w[62][6] ),
    .S0(net445),
    .S1(net1093),
    .X(_02645_));
 sky130_fd_sc_hd__mux4_2 _25866_ (.A0(_02642_),
    .A1(_02643_),
    .A2(_02644_),
    .A3(_02645_),
    .S0(net438),
    .S1(net435),
    .X(_02646_));
 sky130_fd_sc_hd__mux2i_4 _25867_ (.A0(_02641_),
    .A1(_02646_),
    .S(net433),
    .Y(_02647_));
 sky130_fd_sc_hd__xnor2_1 _25868_ (.A(_02621_),
    .B(_02647_),
    .Y(_02648_));
 sky130_fd_sc_hd__xnor2_2 _25869_ (.A(_11451_),
    .B(_02648_),
    .Y(_11736_));
 sky130_fd_sc_hd__xnor2_1 _25870_ (.A(_11220_),
    .B(_11393_),
    .Y(_02649_));
 sky130_fd_sc_hd__xnor2_2 _25871_ (.A(_11104_),
    .B(_02649_),
    .Y(_11739_));
 sky130_fd_sc_hd__mux4_2 _25872_ (.A0(\w[0][7] ),
    .A1(\w[4][7] ),
    .A2(\w[2][7] ),
    .A3(\w[6][7] ),
    .S0(net444),
    .S1(net447),
    .X(_02650_));
 sky130_fd_sc_hd__mux4_2 _25873_ (.A0(\w[8][7] ),
    .A1(\w[12][7] ),
    .A2(\w[10][7] ),
    .A3(\w[14][7] ),
    .S0(net444),
    .S1(net447),
    .X(_02651_));
 sky130_fd_sc_hd__mux4_2 _25874_ (.A0(\w[16][7] ),
    .A1(\w[20][7] ),
    .A2(\w[18][7] ),
    .A3(\w[22][7] ),
    .S0(net444),
    .S1(net447),
    .X(_02652_));
 sky130_fd_sc_hd__mux4_2 _25875_ (.A0(\w[24][7] ),
    .A1(\w[28][7] ),
    .A2(\w[26][7] ),
    .A3(\w[30][7] ),
    .S0(net444),
    .S1(net447),
    .X(_02653_));
 sky130_fd_sc_hd__mux4_2 _25876_ (.A0(_02650_),
    .A1(_02651_),
    .A2(_02652_),
    .A3(_02653_),
    .S0(net437),
    .S1(net435),
    .X(_02654_));
 sky130_fd_sc_hd__mux4_2 _25877_ (.A0(\w[32][7] ),
    .A1(\w[36][7] ),
    .A2(\w[34][7] ),
    .A3(\w[38][7] ),
    .S0(net446),
    .S1(net1093),
    .X(_02655_));
 sky130_fd_sc_hd__mux4_2 _25878_ (.A0(\w[40][7] ),
    .A1(\w[44][7] ),
    .A2(\w[42][7] ),
    .A3(\w[46][7] ),
    .S0(net446),
    .S1(net1093),
    .X(_02656_));
 sky130_fd_sc_hd__mux4_2 _25879_ (.A0(\w[48][7] ),
    .A1(\w[52][7] ),
    .A2(\w[50][7] ),
    .A3(\w[54][7] ),
    .S0(net446),
    .S1(net1093),
    .X(_02657_));
 sky130_fd_sc_hd__mux4_2 _25880_ (.A0(\w[56][7] ),
    .A1(\w[60][7] ),
    .A2(\w[58][7] ),
    .A3(\w[62][7] ),
    .S0(net446),
    .S1(net1093),
    .X(_02658_));
 sky130_fd_sc_hd__mux4_2 _25881_ (.A0(_02655_),
    .A1(_02656_),
    .A2(_02657_),
    .A3(_02658_),
    .S0(net437),
    .S1(net435),
    .X(_02659_));
 sky130_fd_sc_hd__mux2i_4 _25882_ (.A0(_02654_),
    .A1(_02659_),
    .S(net433),
    .Y(_02660_));
 sky130_fd_sc_hd__xnor2_1 _25883_ (.A(_02634_),
    .B(_02660_),
    .Y(_02661_));
 sky130_fd_sc_hd__xnor2_1 _25884_ (.A(_11475_),
    .B(_02661_),
    .Y(_11744_));
 sky130_fd_sc_hd__xnor2_1 _25885_ (.A(_11266_),
    .B(_11439_),
    .Y(_02662_));
 sky130_fd_sc_hd__xnor2_2 _25886_ (.A(_10893_),
    .B(_02662_),
    .Y(_11747_));
 sky130_fd_sc_hd__mux4_2 _25887_ (.A0(\w[0][8] ),
    .A1(\w[4][8] ),
    .A2(\w[2][8] ),
    .A3(\w[6][8] ),
    .S0(net440),
    .S1(net448),
    .X(_02663_));
 sky130_fd_sc_hd__mux4_2 _25888_ (.A0(\w[8][8] ),
    .A1(\w[12][8] ),
    .A2(\w[10][8] ),
    .A3(\w[14][8] ),
    .S0(net440),
    .S1(net448),
    .X(_02664_));
 sky130_fd_sc_hd__mux4_2 _25889_ (.A0(\w[16][8] ),
    .A1(\w[20][8] ),
    .A2(\w[18][8] ),
    .A3(\w[22][8] ),
    .S0(net440),
    .S1(net448),
    .X(_02665_));
 sky130_fd_sc_hd__mux4_2 _25890_ (.A0(\w[24][8] ),
    .A1(\w[28][8] ),
    .A2(\w[26][8] ),
    .A3(\w[30][8] ),
    .S0(net440),
    .S1(net448),
    .X(_02666_));
 sky130_fd_sc_hd__mux4_2 _25891_ (.A0(_02663_),
    .A1(_02664_),
    .A2(_02665_),
    .A3(_02666_),
    .S0(net438),
    .S1(net434),
    .X(_02667_));
 sky130_fd_sc_hd__mux4_2 _25892_ (.A0(\w[32][8] ),
    .A1(\w[36][8] ),
    .A2(\w[34][8] ),
    .A3(\w[38][8] ),
    .S0(net440),
    .S1(net448),
    .X(_02668_));
 sky130_fd_sc_hd__mux4_2 _25893_ (.A0(\w[40][8] ),
    .A1(\w[44][8] ),
    .A2(\w[42][8] ),
    .A3(\w[46][8] ),
    .S0(net440),
    .S1(net448),
    .X(_02669_));
 sky130_fd_sc_hd__mux4_2 _25894_ (.A0(\w[48][8] ),
    .A1(\w[52][8] ),
    .A2(\w[50][8] ),
    .A3(\w[54][8] ),
    .S0(net440),
    .S1(net448),
    .X(_02670_));
 sky130_fd_sc_hd__mux4_2 _25895_ (.A0(\w[56][8] ),
    .A1(\w[60][8] ),
    .A2(\w[58][8] ),
    .A3(\w[62][8] ),
    .S0(net441),
    .S1(net449),
    .X(_02671_));
 sky130_fd_sc_hd__mux4_2 _25896_ (.A0(_02668_),
    .A1(_02669_),
    .A2(_02670_),
    .A3(_02671_),
    .S0(net438),
    .S1(net434),
    .X(_02672_));
 sky130_fd_sc_hd__mux2i_4 _25897_ (.A0(_02667_),
    .A1(_02672_),
    .S(net432),
    .Y(_02673_));
 sky130_fd_sc_hd__xnor2_1 _25898_ (.A(_02647_),
    .B(_02673_),
    .Y(_02674_));
 sky130_fd_sc_hd__xnor2_1 _25899_ (.A(_11499_),
    .B(_02674_),
    .Y(_11752_));
 sky130_fd_sc_hd__xnor2_1 _25900_ (.A(_11323_),
    .B(_11463_),
    .Y(_02675_));
 sky130_fd_sc_hd__xnor2_2 _25901_ (.A(_10917_),
    .B(_02675_),
    .Y(_11755_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_269 ();
 sky130_fd_sc_hd__mux4_2 _25903_ (.A0(\w[0][9] ),
    .A1(\w[4][9] ),
    .A2(\w[2][9] ),
    .A3(\w[6][9] ),
    .S0(net439),
    .S1(net448),
    .X(_02677_));
 sky130_fd_sc_hd__mux4_2 _25904_ (.A0(\w[8][9] ),
    .A1(\w[12][9] ),
    .A2(\w[10][9] ),
    .A3(\w[14][9] ),
    .S0(net439),
    .S1(net448),
    .X(_02678_));
 sky130_fd_sc_hd__mux4_2 _25905_ (.A0(\w[16][9] ),
    .A1(\w[20][9] ),
    .A2(\w[18][9] ),
    .A3(\w[22][9] ),
    .S0(net439),
    .S1(net448),
    .X(_02679_));
 sky130_fd_sc_hd__mux4_2 _25906_ (.A0(\w[24][9] ),
    .A1(\w[28][9] ),
    .A2(\w[26][9] ),
    .A3(\w[30][9] ),
    .S0(net439),
    .S1(net448),
    .X(_02680_));
 sky130_fd_sc_hd__mux4_2 _25907_ (.A0(_02677_),
    .A1(_02678_),
    .A2(_02679_),
    .A3(_02680_),
    .S0(net436),
    .S1(net434),
    .X(_02681_));
 sky130_fd_sc_hd__mux4_2 _25908_ (.A0(\w[32][9] ),
    .A1(\w[36][9] ),
    .A2(\w[34][9] ),
    .A3(\w[38][9] ),
    .S0(net441),
    .S1(net449),
    .X(_02682_));
 sky130_fd_sc_hd__mux4_2 _25909_ (.A0(\w[40][9] ),
    .A1(\w[44][9] ),
    .A2(\w[42][9] ),
    .A3(\w[46][9] ),
    .S0(net441),
    .S1(net449),
    .X(_02683_));
 sky130_fd_sc_hd__mux4_2 _25910_ (.A0(\w[48][9] ),
    .A1(\w[52][9] ),
    .A2(\w[50][9] ),
    .A3(\w[54][9] ),
    .S0(net441),
    .S1(net449),
    .X(_02684_));
 sky130_fd_sc_hd__mux4_2 _25911_ (.A0(\w[56][9] ),
    .A1(\w[60][9] ),
    .A2(\w[58][9] ),
    .A3(\w[62][9] ),
    .S0(net441),
    .S1(net449),
    .X(_02685_));
 sky130_fd_sc_hd__mux4_2 _25912_ (.A0(_02682_),
    .A1(_02683_),
    .A2(_02684_),
    .A3(_02685_),
    .S0(net436),
    .S1(net434),
    .X(_02686_));
 sky130_fd_sc_hd__mux2i_4 _25913_ (.A0(_02681_),
    .A1(_02686_),
    .S(net432),
    .Y(_02687_));
 sky130_fd_sc_hd__xnor2_1 _25914_ (.A(_02660_),
    .B(_02687_),
    .Y(_11760_));
 sky130_fd_sc_hd__xnor2_1 _25915_ (.A(_11358_),
    .B(_11487_),
    .Y(_02688_));
 sky130_fd_sc_hd__xnor2_1 _25916_ (.A(_11045_),
    .B(_02688_),
    .Y(_11763_));
 sky130_fd_sc_hd__mux4_2 _25917_ (.A0(\w[0][10] ),
    .A1(\w[4][10] ),
    .A2(\w[2][10] ),
    .A3(\w[6][10] ),
    .S0(net439),
    .S1(net448),
    .X(_02689_));
 sky130_fd_sc_hd__mux4_2 _25918_ (.A0(\w[8][10] ),
    .A1(\w[12][10] ),
    .A2(\w[10][10] ),
    .A3(\w[14][10] ),
    .S0(net439),
    .S1(net448),
    .X(_02690_));
 sky130_fd_sc_hd__mux4_2 _25919_ (.A0(\w[16][10] ),
    .A1(\w[20][10] ),
    .A2(\w[18][10] ),
    .A3(\w[22][10] ),
    .S0(net439),
    .S1(net448),
    .X(_02691_));
 sky130_fd_sc_hd__mux4_2 _25920_ (.A0(\w[24][10] ),
    .A1(\w[28][10] ),
    .A2(\w[26][10] ),
    .A3(\w[30][10] ),
    .S0(net439),
    .S1(net448),
    .X(_02692_));
 sky130_fd_sc_hd__mux4_2 _25921_ (.A0(_02689_),
    .A1(_02690_),
    .A2(_02691_),
    .A3(_02692_),
    .S0(net436),
    .S1(net434),
    .X(_02693_));
 sky130_fd_sc_hd__mux4_2 _25922_ (.A0(\w[32][10] ),
    .A1(\w[36][10] ),
    .A2(\w[34][10] ),
    .A3(\w[38][10] ),
    .S0(net441),
    .S1(net449),
    .X(_02694_));
 sky130_fd_sc_hd__mux4_2 _25923_ (.A0(\w[40][10] ),
    .A1(\w[44][10] ),
    .A2(\w[42][10] ),
    .A3(\w[46][10] ),
    .S0(net441),
    .S1(net449),
    .X(_02695_));
 sky130_fd_sc_hd__mux4_2 _25924_ (.A0(\w[48][10] ),
    .A1(\w[52][10] ),
    .A2(\w[50][10] ),
    .A3(\w[54][10] ),
    .S0(net441),
    .S1(net449),
    .X(_02696_));
 sky130_fd_sc_hd__mux4_2 _25925_ (.A0(\w[56][10] ),
    .A1(\w[60][10] ),
    .A2(\w[58][10] ),
    .A3(\w[62][10] ),
    .S0(net441),
    .S1(net449),
    .X(_02697_));
 sky130_fd_sc_hd__mux4_2 _25926_ (.A0(_02694_),
    .A1(_02695_),
    .A2(_02696_),
    .A3(_02697_),
    .S0(net436),
    .S1(net434),
    .X(_02698_));
 sky130_fd_sc_hd__mux2i_4 _25927_ (.A0(_02693_),
    .A1(_02698_),
    .S(net432),
    .Y(_02699_));
 sky130_fd_sc_hd__xnor2_1 _25928_ (.A(_02673_),
    .B(_02699_),
    .Y(_11768_));
 sky130_fd_sc_hd__xnor2_1 _25929_ (.A(_11393_),
    .B(_11511_),
    .Y(_02700_));
 sky130_fd_sc_hd__xnor2_2 _25930_ (.A(_11129_),
    .B(_02700_),
    .Y(_11771_));
 sky130_fd_sc_hd__xnor2_1 _25931_ (.A(_10963_),
    .B(_02687_),
    .Y(_11776_));
 sky130_fd_sc_hd__xnor2_1 _25932_ (.A(_11439_),
    .B(_11553_),
    .Y(_02701_));
 sky130_fd_sc_hd__xnor2_2 _25933_ (.A(_11184_),
    .B(_02701_),
    .Y(_11779_));
 sky130_fd_sc_hd__xnor2_1 _25934_ (.A(_11057_),
    .B(_02699_),
    .Y(_11784_));
 sky130_fd_sc_hd__xnor2_1 _25935_ (.A(_11463_),
    .B(_02572_),
    .Y(_02702_));
 sky130_fd_sc_hd__xnor2_1 _25936_ (.A(_11231_),
    .B(_02702_),
    .Y(_11787_));
 sky130_fd_sc_hd__xnor2_1 _25937_ (.A(_10963_),
    .B(_11147_),
    .Y(_11792_));
 sky130_fd_sc_hd__xnor2_1 _25938_ (.A(_11487_),
    .B(_02596_),
    .Y(_02703_));
 sky130_fd_sc_hd__xnor2_1 _25939_ (.A(_11277_),
    .B(_02703_),
    .Y(_11795_));
 sky130_fd_sc_hd__xnor2_1 _25940_ (.A(_11057_),
    .B(_11196_),
    .Y(_11800_));
 sky130_fd_sc_hd__xnor2_1 _25941_ (.A(_11312_),
    .B(_11511_),
    .Y(_02704_));
 sky130_fd_sc_hd__xnor2_1 _25942_ (.A(_10833_),
    .B(_02704_),
    .Y(_11803_));
 sky130_fd_sc_hd__xnor2_1 _25943_ (.A(_11147_),
    .B(_11243_),
    .Y(_11808_));
 sky130_fd_sc_hd__xnor2_1 _25944_ (.A(_10905_),
    .B(_11369_),
    .Y(_11811_));
 sky130_fd_sc_hd__xnor2_1 _25945_ (.A(_11196_),
    .B(_11300_),
    .Y(_11816_));
 sky130_fd_sc_hd__xnor2_1 _25946_ (.A(_11034_),
    .B(_11404_),
    .Y(_11819_));
 sky130_fd_sc_hd__xnor2_1 _25947_ (.A(_11243_),
    .B(_11335_),
    .Y(_11824_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_260 ();
 sky130_fd_sc_hd__mux4_2 _25957_ (.A0(\w[1][10] ),
    .A1(\w[5][10] ),
    .A2(\w[3][10] ),
    .A3(\w[7][10] ),
    .S0(net419),
    .S1(net426),
    .X(_02714_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_258 ();
 sky130_fd_sc_hd__mux4_2 _25960_ (.A0(\w[9][10] ),
    .A1(\w[13][10] ),
    .A2(\w[11][10] ),
    .A3(\w[15][10] ),
    .S0(net419),
    .S1(net426),
    .X(_02717_));
 sky130_fd_sc_hd__mux4_2 _25961_ (.A0(\w[17][10] ),
    .A1(\w[21][10] ),
    .A2(\w[19][10] ),
    .A3(\w[23][10] ),
    .S0(net419),
    .S1(net426),
    .X(_02718_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_255 ();
 sky130_fd_sc_hd__mux4_2 _25965_ (.A0(\w[25][10] ),
    .A1(\w[29][10] ),
    .A2(\w[27][10] ),
    .A3(\w[31][10] ),
    .S0(net419),
    .S1(net426),
    .X(_02722_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_250 ();
 sky130_fd_sc_hd__mux4_2 _25971_ (.A0(_02714_),
    .A1(_02717_),
    .A2(_02718_),
    .A3(_02722_),
    .S0(net418),
    .S1(net415),
    .X(_02728_));
 sky130_fd_sc_hd__mux4_2 _25972_ (.A0(\w[33][10] ),
    .A1(\w[37][10] ),
    .A2(\w[35][10] ),
    .A3(\w[39][10] ),
    .S0(net421),
    .S1(net428),
    .X(_02729_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_248 ();
 sky130_fd_sc_hd__mux4_2 _25975_ (.A0(\w[41][10] ),
    .A1(\w[45][10] ),
    .A2(\w[43][10] ),
    .A3(\w[47][10] ),
    .S0(net421),
    .S1(net428),
    .X(_02732_));
 sky130_fd_sc_hd__mux4_2 _25976_ (.A0(\w[49][10] ),
    .A1(\w[53][10] ),
    .A2(\w[51][10] ),
    .A3(\w[55][10] ),
    .S0(net421),
    .S1(net428),
    .X(_02733_));
 sky130_fd_sc_hd__mux4_2 _25977_ (.A0(\w[57][10] ),
    .A1(\w[61][10] ),
    .A2(\w[59][10] ),
    .A3(\w[63][10] ),
    .S0(net421),
    .S1(net428),
    .X(_02734_));
 sky130_fd_sc_hd__mux4_2 _25978_ (.A0(_02729_),
    .A1(_02732_),
    .A2(_02733_),
    .A3(_02734_),
    .S0(net418),
    .S1(net415),
    .X(_02735_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_246 ();
 sky130_fd_sc_hd__mux2i_4 _25981_ (.A0(_02728_),
    .A1(_02735_),
    .S(net539),
    .Y(_02738_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_243 ();
 sky130_fd_sc_hd__mux4_2 _25985_ (.A0(\w[1][19] ),
    .A1(\w[5][19] ),
    .A2(\w[3][19] ),
    .A3(\w[7][19] ),
    .S0(net419),
    .S1(net426),
    .X(_02742_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_241 ();
 sky130_fd_sc_hd__mux4_2 _25988_ (.A0(\w[9][19] ),
    .A1(\w[13][19] ),
    .A2(\w[11][19] ),
    .A3(\w[15][19] ),
    .S0(net419),
    .S1(net426),
    .X(_02745_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_239 ();
 sky130_fd_sc_hd__mux4_2 _25991_ (.A0(\w[17][19] ),
    .A1(\w[21][19] ),
    .A2(\w[19][19] ),
    .A3(\w[23][19] ),
    .S0(net419),
    .S1(net426),
    .X(_02748_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_237 ();
 sky130_fd_sc_hd__mux4_2 _25994_ (.A0(\w[25][19] ),
    .A1(\w[29][19] ),
    .A2(\w[27][19] ),
    .A3(\w[31][19] ),
    .S0(net419),
    .S1(net426),
    .X(_02751_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_235 ();
 sky130_fd_sc_hd__mux4_2 _25997_ (.A0(_02742_),
    .A1(_02745_),
    .A2(_02748_),
    .A3(_02751_),
    .S0(net418),
    .S1(net415),
    .X(_02754_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_234 ();
 sky130_fd_sc_hd__mux4_2 _25999_ (.A0(\w[33][19] ),
    .A1(\w[37][19] ),
    .A2(\w[35][19] ),
    .A3(\w[39][19] ),
    .S0(net421),
    .S1(net428),
    .X(_02756_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_232 ();
 sky130_fd_sc_hd__mux4_2 _26002_ (.A0(\w[41][19] ),
    .A1(\w[45][19] ),
    .A2(\w[43][19] ),
    .A3(\w[47][19] ),
    .S0(net421),
    .S1(net428),
    .X(_02759_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_230 ();
 sky130_fd_sc_hd__mux4_2 _26005_ (.A0(\w[49][19] ),
    .A1(\w[53][19] ),
    .A2(\w[51][19] ),
    .A3(\w[55][19] ),
    .S0(net421),
    .S1(net428),
    .X(_02762_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_228 ();
 sky130_fd_sc_hd__mux4_2 _26008_ (.A0(\w[57][19] ),
    .A1(\w[61][19] ),
    .A2(\w[59][19] ),
    .A3(\w[63][19] ),
    .S0(net421),
    .S1(net428),
    .X(_02765_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_226 ();
 sky130_fd_sc_hd__mux4_2 _26011_ (.A0(_02756_),
    .A1(_02759_),
    .A2(_02762_),
    .A3(_02765_),
    .S0(net418),
    .S1(net415),
    .X(_02768_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_225 ();
 sky130_fd_sc_hd__mux2i_4 _26013_ (.A0(_02754_),
    .A1(_02768_),
    .S(net539),
    .Y(_02770_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_224 ();
 sky130_fd_sc_hd__mux4_2 _26015_ (.A0(\w[1][17] ),
    .A1(\w[5][17] ),
    .A2(\w[3][17] ),
    .A3(\w[7][17] ),
    .S0(net422),
    .S1(net429),
    .X(_02772_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_222 ();
 sky130_fd_sc_hd__mux4_2 _26018_ (.A0(\w[9][17] ),
    .A1(\w[13][17] ),
    .A2(\w[11][17] ),
    .A3(\w[15][17] ),
    .S0(net422),
    .S1(net429),
    .X(_02775_));
 sky130_fd_sc_hd__mux4_2 _26019_ (.A0(\w[17][17] ),
    .A1(\w[21][17] ),
    .A2(\w[19][17] ),
    .A3(\w[23][17] ),
    .S0(net422),
    .S1(net429),
    .X(_02776_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_220 ();
 sky130_fd_sc_hd__mux4_2 _26022_ (.A0(\w[25][17] ),
    .A1(\w[29][17] ),
    .A2(\w[27][17] ),
    .A3(\w[31][17] ),
    .S0(net422),
    .S1(net429),
    .X(_02779_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_218 ();
 sky130_fd_sc_hd__mux4_2 _26025_ (.A0(_02772_),
    .A1(_02775_),
    .A2(_02776_),
    .A3(_02779_),
    .S0(net416),
    .S1(net414),
    .X(_02782_));
 sky130_fd_sc_hd__mux4_2 _26026_ (.A0(\w[33][17] ),
    .A1(\w[37][17] ),
    .A2(\w[35][17] ),
    .A3(\w[39][17] ),
    .S0(net422),
    .S1(net429),
    .X(_02783_));
 sky130_fd_sc_hd__mux4_2 _26027_ (.A0(\w[41][17] ),
    .A1(\w[45][17] ),
    .A2(\w[43][17] ),
    .A3(\w[47][17] ),
    .S0(net422),
    .S1(net429),
    .X(_02784_));
 sky130_fd_sc_hd__mux4_2 _26028_ (.A0(\w[49][17] ),
    .A1(\w[53][17] ),
    .A2(\w[51][17] ),
    .A3(\w[55][17] ),
    .S0(net422),
    .S1(net429),
    .X(_02785_));
 sky130_fd_sc_hd__mux4_2 _26029_ (.A0(\w[57][17] ),
    .A1(\w[61][17] ),
    .A2(\w[59][17] ),
    .A3(\w[63][17] ),
    .S0(net422),
    .S1(net429),
    .X(_02786_));
 sky130_fd_sc_hd__mux4_2 _26030_ (.A0(_02783_),
    .A1(_02784_),
    .A2(_02785_),
    .A3(_02786_),
    .S0(net416),
    .S1(net414),
    .X(_02787_));
 sky130_fd_sc_hd__mux2i_4 _26031_ (.A0(_02782_),
    .A1(_02787_),
    .S(net413),
    .Y(_02788_));
 sky130_fd_sc_hd__xnor2_1 _26032_ (.A(_02770_),
    .B(_02788_),
    .Y(_02789_));
 sky130_fd_sc_hd__xnor2_1 _26033_ (.A(_02738_),
    .B(_02789_),
    .Y(_11829_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_209 ();
 sky130_fd_sc_hd__mux4_2 _26043_ (.A0(\w[0][3] ),
    .A1(\w[4][3] ),
    .A2(\w[2][3] ),
    .A3(\w[6][3] ),
    .S0(net1133),
    .S1(\count15_2[1] ),
    .X(_02799_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_205 ();
 sky130_fd_sc_hd__mux4_2 _26048_ (.A0(\w[8][3] ),
    .A1(\w[12][3] ),
    .A2(\w[10][3] ),
    .A3(\w[14][3] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_02804_));
 sky130_fd_sc_hd__mux4_2 _26049_ (.A0(\w[16][3] ),
    .A1(\w[20][3] ),
    .A2(\w[18][3] ),
    .A3(\w[22][3] ),
    .S0(net1133),
    .S1(\count15_2[1] ),
    .X(_02805_));
 sky130_fd_sc_hd__mux4_2 _26050_ (.A0(\w[24][3] ),
    .A1(\w[28][3] ),
    .A2(\w[26][3] ),
    .A3(\w[30][3] ),
    .S0(\count15_2[2] ),
    .S1(\count15_2[1] ),
    .X(_02806_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_200 ();
 sky130_fd_sc_hd__mux4_2 _26056_ (.A0(_02799_),
    .A1(_02804_),
    .A2(_02805_),
    .A3(_02806_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[4] ),
    .X(_02812_));
 sky130_fd_sc_hd__mux4_2 _26057_ (.A0(\w[32][3] ),
    .A1(\w[36][3] ),
    .A2(\w[34][3] ),
    .A3(\w[38][3] ),
    .S0(net505),
    .S1(\count15_2[1] ),
    .X(_02813_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_196 ();
 sky130_fd_sc_hd__mux4_2 _26062_ (.A0(\w[40][3] ),
    .A1(\w[44][3] ),
    .A2(\w[42][3] ),
    .A3(\w[46][3] ),
    .S0(net505),
    .S1(\count15_2[1] ),
    .X(_02818_));
 sky130_fd_sc_hd__mux4_2 _26063_ (.A0(\w[48][3] ),
    .A1(\w[52][3] ),
    .A2(\w[50][3] ),
    .A3(\w[54][3] ),
    .S0(net505),
    .S1(\count15_2[1] ),
    .X(_02819_));
 sky130_fd_sc_hd__mux4_2 _26064_ (.A0(\w[56][3] ),
    .A1(\w[60][3] ),
    .A2(\w[58][3] ),
    .A3(\w[62][3] ),
    .S0(net505),
    .S1(\count15_2[1] ),
    .X(_02820_));
 sky130_fd_sc_hd__mux4_2 _26065_ (.A0(_02813_),
    .A1(_02818_),
    .A2(_02819_),
    .A3(_02820_),
    .S0(net497),
    .S1(\count15_2[4] ),
    .X(_02821_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_194 ();
 sky130_fd_sc_hd__mux2i_4 _26068_ (.A0(_02812_),
    .A1(_02821_),
    .S(\count15_2[5] ),
    .Y(_02824_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_192 ();
 sky130_fd_sc_hd__mux4_2 _26071_ (.A0(\w[0][18] ),
    .A1(\w[4][18] ),
    .A2(\w[2][18] ),
    .A3(\w[6][18] ),
    .S0(net504),
    .S1(net510),
    .X(_02827_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_190 ();
 sky130_fd_sc_hd__mux4_2 _26074_ (.A0(\w[8][18] ),
    .A1(\w[12][18] ),
    .A2(\w[10][18] ),
    .A3(\w[14][18] ),
    .S0(net504),
    .S1(net510),
    .X(_02830_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_188 ();
 sky130_fd_sc_hd__mux4_2 _26077_ (.A0(\w[16][18] ),
    .A1(\w[20][18] ),
    .A2(\w[18][18] ),
    .A3(\w[22][18] ),
    .S0(net504),
    .S1(net510),
    .X(_02833_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_186 ();
 sky130_fd_sc_hd__mux4_2 _26080_ (.A0(\w[24][18] ),
    .A1(\w[28][18] ),
    .A2(\w[26][18] ),
    .A3(\w[30][18] ),
    .S0(net504),
    .S1(net510),
    .X(_02836_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_184 ();
 sky130_fd_sc_hd__mux4_2 _26083_ (.A0(_02827_),
    .A1(_02830_),
    .A2(_02833_),
    .A3(_02836_),
    .S0(net497),
    .S1(net495),
    .X(_02839_));
 sky130_fd_sc_hd__mux4_2 _26084_ (.A0(\w[32][18] ),
    .A1(\w[36][18] ),
    .A2(\w[34][18] ),
    .A3(\w[38][18] ),
    .S0(net504),
    .S1(net510),
    .X(_02840_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_183 ();
 sky130_fd_sc_hd__mux4_2 _26086_ (.A0(\w[40][18] ),
    .A1(\w[44][18] ),
    .A2(\w[42][18] ),
    .A3(\w[46][18] ),
    .S0(net504),
    .S1(net510),
    .X(_02842_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_181 ();
 sky130_fd_sc_hd__mux4_2 _26089_ (.A0(\w[48][18] ),
    .A1(\w[52][18] ),
    .A2(\w[50][18] ),
    .A3(\w[54][18] ),
    .S0(net504),
    .S1(net510),
    .X(_02845_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_179 ();
 sky130_fd_sc_hd__mux4_2 _26092_ (.A0(\w[56][18] ),
    .A1(\w[60][18] ),
    .A2(\w[58][18] ),
    .A3(\w[62][18] ),
    .S0(net504),
    .S1(net510),
    .X(_02848_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_177 ();
 sky130_fd_sc_hd__mux4_2 _26095_ (.A0(_02840_),
    .A1(_02842_),
    .A2(_02845_),
    .A3(_02848_),
    .S0(net497),
    .S1(net495),
    .X(_02851_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_176 ();
 sky130_fd_sc_hd__mux2i_4 _26097_ (.A0(_02839_),
    .A1(_02851_),
    .S(net492),
    .Y(_02853_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_174 ();
 sky130_fd_sc_hd__mux4_2 _26100_ (.A0(\w[0][7] ),
    .A1(\w[4][7] ),
    .A2(\w[2][7] ),
    .A3(\w[6][7] ),
    .S0(net498),
    .S1(net506),
    .X(_02856_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_172 ();
 sky130_fd_sc_hd__mux4_2 _26103_ (.A0(\w[8][7] ),
    .A1(\w[12][7] ),
    .A2(\w[10][7] ),
    .A3(\w[14][7] ),
    .S0(net499),
    .S1(net506),
    .X(_02859_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_171 ();
 sky130_fd_sc_hd__mux4_2 _26105_ (.A0(\w[16][7] ),
    .A1(\w[20][7] ),
    .A2(\w[18][7] ),
    .A3(\w[22][7] ),
    .S0(net498),
    .S1(net506),
    .X(_02861_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_170 ();
 sky130_fd_sc_hd__mux4_2 _26107_ (.A0(\w[24][7] ),
    .A1(\w[28][7] ),
    .A2(\w[26][7] ),
    .A3(\w[30][7] ),
    .S0(net499),
    .S1(net506),
    .X(_02863_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_168 ();
 sky130_fd_sc_hd__mux4_2 _26110_ (.A0(_02856_),
    .A1(_02859_),
    .A2(_02861_),
    .A3(_02863_),
    .S0(net496),
    .S1(net547),
    .X(_02866_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_166 ();
 sky130_fd_sc_hd__mux4_2 _26113_ (.A0(\w[32][7] ),
    .A1(\w[36][7] ),
    .A2(\w[34][7] ),
    .A3(\w[38][7] ),
    .S0(net505),
    .S1(\count15_2[1] ),
    .X(_02869_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_164 ();
 sky130_fd_sc_hd__mux4_2 _26116_ (.A0(\w[40][7] ),
    .A1(\w[44][7] ),
    .A2(\w[42][7] ),
    .A3(\w[46][7] ),
    .S0(net505),
    .S1(\count15_2[1] ),
    .X(_02872_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_162 ();
 sky130_fd_sc_hd__mux4_2 _26119_ (.A0(\w[48][7] ),
    .A1(\w[52][7] ),
    .A2(\w[50][7] ),
    .A3(\w[54][7] ),
    .S0(net505),
    .S1(\count15_2[1] ),
    .X(_02875_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_160 ();
 sky130_fd_sc_hd__mux4_2 _26122_ (.A0(\w[56][7] ),
    .A1(\w[60][7] ),
    .A2(\w[58][7] ),
    .A3(\w[62][7] ),
    .S0(net505),
    .S1(\count15_2[1] ),
    .X(_02878_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_158 ();
 sky130_fd_sc_hd__mux4_2 _26125_ (.A0(_02869_),
    .A1(_02872_),
    .A2(_02875_),
    .A3(_02878_),
    .S0(\count15_2[3] ),
    .S1(net547),
    .X(_02881_));
 sky130_fd_sc_hd__mux2i_4 _26126_ (.A0(_02866_),
    .A1(_02881_),
    .S(net493),
    .Y(_02882_));
 sky130_fd_sc_hd__xnor2_1 _26127_ (.A(_02853_),
    .B(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__xnor2_2 _26128_ (.A(_02824_),
    .B(_02883_),
    .Y(_11828_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_150 ();
 sky130_fd_sc_hd__mux4_2 _26137_ (.A0(\w[0][0] ),
    .A1(\w[4][0] ),
    .A2(\w[2][0] ),
    .A3(\w[6][0] ),
    .S0(net381),
    .S1(net389),
    .X(_02892_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_146 ();
 sky130_fd_sc_hd__mux4_2 _26142_ (.A0(\w[8][0] ),
    .A1(\w[12][0] ),
    .A2(\w[10][0] ),
    .A3(\w[14][0] ),
    .S0(net381),
    .S1(net389),
    .X(_02897_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_144 ();
 sky130_fd_sc_hd__mux4_2 _26145_ (.A0(\w[16][0] ),
    .A1(\w[20][0] ),
    .A2(\w[18][0] ),
    .A3(\w[22][0] ),
    .S0(net381),
    .S1(net389),
    .X(_02900_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_141 ();
 sky130_fd_sc_hd__mux4_2 _26149_ (.A0(\w[24][0] ),
    .A1(\w[28][0] ),
    .A2(\w[26][0] ),
    .A3(\w[30][0] ),
    .S0(net381),
    .S1(net389),
    .X(_02904_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_136 ();
 sky130_fd_sc_hd__mux4_2 _26155_ (.A0(_02892_),
    .A1(_02897_),
    .A2(_02900_),
    .A3(_02904_),
    .S0(net378),
    .S1(net535),
    .X(_02910_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_134 ();
 sky130_fd_sc_hd__mux4_2 _26158_ (.A0(\w[32][0] ),
    .A1(\w[36][0] ),
    .A2(\w[34][0] ),
    .A3(\w[38][0] ),
    .S0(net383),
    .S1(net390),
    .X(_02913_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_132 ();
 sky130_fd_sc_hd__mux4_2 _26161_ (.A0(\w[40][0] ),
    .A1(\w[44][0] ),
    .A2(\w[42][0] ),
    .A3(\w[46][0] ),
    .S0(net383),
    .S1(net390),
    .X(_02916_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_130 ();
 sky130_fd_sc_hd__mux4_2 _26164_ (.A0(\w[48][0] ),
    .A1(\w[52][0] ),
    .A2(\w[50][0] ),
    .A3(\w[54][0] ),
    .S0(net383),
    .S1(net390),
    .X(_02919_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_128 ();
 sky130_fd_sc_hd__mux4_2 _26167_ (.A0(\w[56][0] ),
    .A1(\w[60][0] ),
    .A2(\w[58][0] ),
    .A3(\w[62][0] ),
    .S0(net383),
    .S1(net390),
    .X(_02922_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_126 ();
 sky130_fd_sc_hd__mux4_2 _26170_ (.A0(_02913_),
    .A1(_02916_),
    .A2(_02919_),
    .A3(_02922_),
    .S0(net378),
    .S1(net535),
    .X(_02925_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_124 ();
 sky130_fd_sc_hd__mux2i_4 _26173_ (.A0(_02910_),
    .A1(_02925_),
    .S(net374),
    .Y(_11827_));
 sky130_fd_sc_hd__mux4_2 _26174_ (.A0(\w[1][11] ),
    .A1(\w[5][11] ),
    .A2(\w[3][11] ),
    .A3(\w[7][11] ),
    .S0(net420),
    .S1(net427),
    .X(_02928_));
 sky130_fd_sc_hd__mux4_2 _26175_ (.A0(\w[9][11] ),
    .A1(\w[13][11] ),
    .A2(\w[11][11] ),
    .A3(\w[15][11] ),
    .S0(net420),
    .S1(net427),
    .X(_02929_));
 sky130_fd_sc_hd__mux4_2 _26176_ (.A0(\w[17][11] ),
    .A1(\w[21][11] ),
    .A2(\w[19][11] ),
    .A3(\w[23][11] ),
    .S0(net420),
    .S1(net427),
    .X(_02930_));
 sky130_fd_sc_hd__mux4_2 _26177_ (.A0(\w[25][11] ),
    .A1(\w[29][11] ),
    .A2(\w[27][11] ),
    .A3(\w[31][11] ),
    .S0(net420),
    .S1(net427),
    .X(_02931_));
 sky130_fd_sc_hd__mux4_2 _26178_ (.A0(_02928_),
    .A1(_02929_),
    .A2(_02930_),
    .A3(_02931_),
    .S0(net416),
    .S1(net415),
    .X(_02932_));
 sky130_fd_sc_hd__mux4_2 _26179_ (.A0(\w[33][11] ),
    .A1(\w[37][11] ),
    .A2(\w[35][11] ),
    .A3(\w[39][11] ),
    .S0(net425),
    .S1(net430),
    .X(_02933_));
 sky130_fd_sc_hd__mux4_2 _26180_ (.A0(\w[41][11] ),
    .A1(\w[45][11] ),
    .A2(\w[43][11] ),
    .A3(\w[47][11] ),
    .S0(net425),
    .S1(net430),
    .X(_02934_));
 sky130_fd_sc_hd__mux4_2 _26181_ (.A0(\w[49][11] ),
    .A1(\w[53][11] ),
    .A2(\w[51][11] ),
    .A3(\w[55][11] ),
    .S0(net425),
    .S1(net430),
    .X(_02935_));
 sky130_fd_sc_hd__mux4_2 _26182_ (.A0(\w[57][11] ),
    .A1(\w[61][11] ),
    .A2(\w[59][11] ),
    .A3(\w[63][11] ),
    .S0(net425),
    .S1(net430),
    .X(_02936_));
 sky130_fd_sc_hd__mux4_2 _26183_ (.A0(_02933_),
    .A1(_02934_),
    .A2(_02935_),
    .A3(_02936_),
    .S0(net418),
    .S1(net415),
    .X(_02937_));
 sky130_fd_sc_hd__mux2i_4 _26184_ (.A0(_02932_),
    .A1(_02937_),
    .S(net539),
    .Y(_02938_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_123 ();
 sky130_fd_sc_hd__mux4_2 _26186_ (.A0(\w[1][20] ),
    .A1(\w[5][20] ),
    .A2(\w[3][20] ),
    .A3(\w[7][20] ),
    .S0(net421),
    .S1(net428),
    .X(_02940_));
 sky130_fd_sc_hd__mux4_2 _26187_ (.A0(\w[9][20] ),
    .A1(\w[13][20] ),
    .A2(\w[11][20] ),
    .A3(\w[15][20] ),
    .S0(net421),
    .S1(net428),
    .X(_02941_));
 sky130_fd_sc_hd__mux4_2 _26188_ (.A0(\w[17][20] ),
    .A1(\w[21][20] ),
    .A2(\w[19][20] ),
    .A3(\w[23][20] ),
    .S0(net421),
    .S1(net428),
    .X(_02942_));
 sky130_fd_sc_hd__mux4_2 _26189_ (.A0(\w[25][20] ),
    .A1(\w[29][20] ),
    .A2(\w[27][20] ),
    .A3(\w[31][20] ),
    .S0(net421),
    .S1(net428),
    .X(_02943_));
 sky130_fd_sc_hd__mux4_2 _26190_ (.A0(_02940_),
    .A1(_02941_),
    .A2(_02942_),
    .A3(_02943_),
    .S0(net418),
    .S1(net415),
    .X(_02944_));
 sky130_fd_sc_hd__mux4_2 _26191_ (.A0(\w[33][20] ),
    .A1(\w[37][20] ),
    .A2(\w[35][20] ),
    .A3(\w[39][20] ),
    .S0(net425),
    .S1(net430),
    .X(_02945_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_122 ();
 sky130_fd_sc_hd__mux4_2 _26193_ (.A0(\w[41][20] ),
    .A1(\w[45][20] ),
    .A2(\w[43][20] ),
    .A3(\w[47][20] ),
    .S0(net425),
    .S1(net430),
    .X(_02947_));
 sky130_fd_sc_hd__mux4_2 _26194_ (.A0(\w[49][20] ),
    .A1(\w[53][20] ),
    .A2(\w[51][20] ),
    .A3(\w[55][20] ),
    .S0(net425),
    .S1(net430),
    .X(_02948_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_121 ();
 sky130_fd_sc_hd__mux4_2 _26196_ (.A0(\w[57][20] ),
    .A1(\w[61][20] ),
    .A2(\w[59][20] ),
    .A3(\w[63][20] ),
    .S0(net425),
    .S1(net430),
    .X(_02950_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_120 ();
 sky130_fd_sc_hd__mux4_2 _26198_ (.A0(_02945_),
    .A1(_02947_),
    .A2(_02948_),
    .A3(_02950_),
    .S0(net418),
    .S1(net415),
    .X(_02952_));
 sky130_fd_sc_hd__mux2i_4 _26199_ (.A0(_02944_),
    .A1(_02952_),
    .S(net539),
    .Y(_02953_));
 sky130_fd_sc_hd__mux4_2 _26200_ (.A0(\w[1][18] ),
    .A1(\w[5][18] ),
    .A2(\w[3][18] ),
    .A3(\w[7][18] ),
    .S0(net419),
    .S1(net426),
    .X(_02954_));
 sky130_fd_sc_hd__mux4_2 _26201_ (.A0(\w[9][18] ),
    .A1(\w[13][18] ),
    .A2(\w[11][18] ),
    .A3(\w[15][18] ),
    .S0(net419),
    .S1(net426),
    .X(_02955_));
 sky130_fd_sc_hd__mux4_2 _26202_ (.A0(\w[17][18] ),
    .A1(\w[21][18] ),
    .A2(\w[19][18] ),
    .A3(\w[23][18] ),
    .S0(net419),
    .S1(net426),
    .X(_02956_));
 sky130_fd_sc_hd__mux4_2 _26203_ (.A0(\w[25][18] ),
    .A1(\w[29][18] ),
    .A2(\w[27][18] ),
    .A3(\w[31][18] ),
    .S0(net419),
    .S1(net426),
    .X(_02957_));
 sky130_fd_sc_hd__mux4_2 _26204_ (.A0(_02954_),
    .A1(_02955_),
    .A2(_02956_),
    .A3(_02957_),
    .S0(net418),
    .S1(net415),
    .X(_02958_));
 sky130_fd_sc_hd__mux4_2 _26205_ (.A0(\w[33][18] ),
    .A1(\w[37][18] ),
    .A2(\w[35][18] ),
    .A3(\w[39][18] ),
    .S0(net421),
    .S1(net428),
    .X(_02959_));
 sky130_fd_sc_hd__mux4_2 _26206_ (.A0(\w[41][18] ),
    .A1(\w[45][18] ),
    .A2(\w[43][18] ),
    .A3(\w[47][18] ),
    .S0(net421),
    .S1(net428),
    .X(_02960_));
 sky130_fd_sc_hd__mux4_2 _26207_ (.A0(\w[49][18] ),
    .A1(\w[53][18] ),
    .A2(\w[51][18] ),
    .A3(\w[55][18] ),
    .S0(net421),
    .S1(net428),
    .X(_02961_));
 sky130_fd_sc_hd__mux4_2 _26208_ (.A0(\w[57][18] ),
    .A1(\w[61][18] ),
    .A2(\w[59][18] ),
    .A3(\w[63][18] ),
    .S0(net421),
    .S1(net428),
    .X(_02962_));
 sky130_fd_sc_hd__mux4_2 _26209_ (.A0(_02959_),
    .A1(_02960_),
    .A2(_02961_),
    .A3(_02962_),
    .S0(net418),
    .S1(net415),
    .X(_02963_));
 sky130_fd_sc_hd__mux2i_4 _26210_ (.A0(_02958_),
    .A1(_02963_),
    .S(net539),
    .Y(_02964_));
 sky130_fd_sc_hd__xnor2_1 _26211_ (.A(_02953_),
    .B(_02964_),
    .Y(_02965_));
 sky130_fd_sc_hd__xnor2_1 _26212_ (.A(_02938_),
    .B(_02965_),
    .Y(_11834_));
 sky130_fd_sc_hd__mux4_2 _26213_ (.A0(\w[0][4] ),
    .A1(\w[4][4] ),
    .A2(\w[2][4] ),
    .A3(\w[6][4] ),
    .S0(net499),
    .S1(net506),
    .X(_02966_));
 sky130_fd_sc_hd__mux4_2 _26214_ (.A0(\w[8][4] ),
    .A1(\w[12][4] ),
    .A2(\w[10][4] ),
    .A3(\w[14][4] ),
    .S0(net499),
    .S1(net506),
    .X(_02967_));
 sky130_fd_sc_hd__mux4_2 _26215_ (.A0(\w[16][4] ),
    .A1(\w[20][4] ),
    .A2(\w[18][4] ),
    .A3(\w[22][4] ),
    .S0(net499),
    .S1(net506),
    .X(_02968_));
 sky130_fd_sc_hd__mux4_2 _26216_ (.A0(\w[24][4] ),
    .A1(\w[28][4] ),
    .A2(\w[26][4] ),
    .A3(\w[30][4] ),
    .S0(net499),
    .S1(net506),
    .X(_02969_));
 sky130_fd_sc_hd__mux4_2 _26217_ (.A0(_02966_),
    .A1(_02967_),
    .A2(_02968_),
    .A3(_02969_),
    .S0(net496),
    .S1(net547),
    .X(_02970_));
 sky130_fd_sc_hd__mux4_2 _26218_ (.A0(\w[32][4] ),
    .A1(\w[36][4] ),
    .A2(\w[34][4] ),
    .A3(\w[38][4] ),
    .S0(net499),
    .S1(net506),
    .X(_02971_));
 sky130_fd_sc_hd__mux4_2 _26219_ (.A0(\w[40][4] ),
    .A1(\w[44][4] ),
    .A2(\w[42][4] ),
    .A3(\w[46][4] ),
    .S0(net499),
    .S1(net506),
    .X(_02972_));
 sky130_fd_sc_hd__mux4_2 _26220_ (.A0(\w[48][4] ),
    .A1(\w[52][4] ),
    .A2(\w[50][4] ),
    .A3(\w[54][4] ),
    .S0(net499),
    .S1(net506),
    .X(_02973_));
 sky130_fd_sc_hd__mux4_2 _26221_ (.A0(\w[56][4] ),
    .A1(\w[60][4] ),
    .A2(\w[58][4] ),
    .A3(\w[62][4] ),
    .S0(net499),
    .S1(net506),
    .X(_02974_));
 sky130_fd_sc_hd__mux4_2 _26222_ (.A0(_02971_),
    .A1(_02972_),
    .A2(_02973_),
    .A3(_02974_),
    .S0(net496),
    .S1(net547),
    .X(_02975_));
 sky130_fd_sc_hd__mux2i_4 _26223_ (.A0(_02970_),
    .A1(_02975_),
    .S(net493),
    .Y(_02976_));
 sky130_fd_sc_hd__mux4_2 _26224_ (.A0(\w[0][8] ),
    .A1(\w[4][8] ),
    .A2(\w[2][8] ),
    .A3(\w[6][8] ),
    .S0(net501),
    .S1(net507),
    .X(_02977_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_118 ();
 sky130_fd_sc_hd__mux4_2 _26227_ (.A0(\w[8][8] ),
    .A1(\w[12][8] ),
    .A2(\w[10][8] ),
    .A3(\w[14][8] ),
    .S0(net501),
    .S1(net507),
    .X(_02980_));
 sky130_fd_sc_hd__mux4_2 _26228_ (.A0(\w[16][8] ),
    .A1(\w[20][8] ),
    .A2(\w[18][8] ),
    .A3(\w[22][8] ),
    .S0(net501),
    .S1(net507),
    .X(_02981_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_117 ();
 sky130_fd_sc_hd__mux4_2 _26230_ (.A0(\w[24][8] ),
    .A1(\w[28][8] ),
    .A2(\w[26][8] ),
    .A3(\w[30][8] ),
    .S0(net501),
    .S1(net507),
    .X(_02983_));
 sky130_fd_sc_hd__mux4_2 _26231_ (.A0(_02977_),
    .A1(_02980_),
    .A2(_02981_),
    .A3(_02983_),
    .S0(net496),
    .S1(net494),
    .X(_02984_));
 sky130_fd_sc_hd__mux4_2 _26232_ (.A0(\w[32][8] ),
    .A1(\w[36][8] ),
    .A2(\w[34][8] ),
    .A3(\w[38][8] ),
    .S0(net501),
    .S1(net507),
    .X(_02985_));
 sky130_fd_sc_hd__mux4_2 _26233_ (.A0(\w[40][8] ),
    .A1(\w[44][8] ),
    .A2(\w[42][8] ),
    .A3(\w[46][8] ),
    .S0(net501),
    .S1(net507),
    .X(_02986_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_115 ();
 sky130_fd_sc_hd__mux4_2 _26236_ (.A0(\w[48][8] ),
    .A1(\w[52][8] ),
    .A2(\w[50][8] ),
    .A3(\w[54][8] ),
    .S0(net501),
    .S1(net507),
    .X(_02989_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_113 ();
 sky130_fd_sc_hd__mux4_2 _26239_ (.A0(\w[56][8] ),
    .A1(\w[60][8] ),
    .A2(\w[58][8] ),
    .A3(\w[62][8] ),
    .S0(net502),
    .S1(net508),
    .X(_02992_));
 sky130_fd_sc_hd__mux4_2 _26240_ (.A0(_02985_),
    .A1(_02986_),
    .A2(_02989_),
    .A3(_02992_),
    .S0(net548),
    .S1(net494),
    .X(_02993_));
 sky130_fd_sc_hd__mux2i_4 _26241_ (.A0(_02984_),
    .A1(_02993_),
    .S(net492),
    .Y(_02994_));
 sky130_fd_sc_hd__mux4_2 _26242_ (.A0(\w[0][19] ),
    .A1(\w[4][19] ),
    .A2(\w[2][19] ),
    .A3(\w[6][19] ),
    .S0(net501),
    .S1(net507),
    .X(_02995_));
 sky130_fd_sc_hd__mux4_2 _26243_ (.A0(\w[8][19] ),
    .A1(\w[12][19] ),
    .A2(\w[10][19] ),
    .A3(\w[14][19] ),
    .S0(net501),
    .S1(net507),
    .X(_02996_));
 sky130_fd_sc_hd__mux4_2 _26244_ (.A0(\w[16][19] ),
    .A1(\w[20][19] ),
    .A2(\w[18][19] ),
    .A3(\w[22][19] ),
    .S0(net501),
    .S1(net507),
    .X(_02997_));
 sky130_fd_sc_hd__mux4_2 _26245_ (.A0(\w[24][19] ),
    .A1(\w[28][19] ),
    .A2(\w[26][19] ),
    .A3(\w[30][19] ),
    .S0(net501),
    .S1(net507),
    .X(_02998_));
 sky130_fd_sc_hd__mux4_2 _26246_ (.A0(_02995_),
    .A1(_02996_),
    .A2(_02997_),
    .A3(_02998_),
    .S0(net496),
    .S1(net494),
    .X(_02999_));
 sky130_fd_sc_hd__mux4_2 _26247_ (.A0(\w[32][19] ),
    .A1(\w[36][19] ),
    .A2(\w[34][19] ),
    .A3(\w[38][19] ),
    .S0(net502),
    .S1(net508),
    .X(_03000_));
 sky130_fd_sc_hd__mux4_2 _26248_ (.A0(\w[40][19] ),
    .A1(\w[44][19] ),
    .A2(\w[42][19] ),
    .A3(\w[46][19] ),
    .S0(net502),
    .S1(net508),
    .X(_03001_));
 sky130_fd_sc_hd__mux4_2 _26249_ (.A0(\w[48][19] ),
    .A1(\w[52][19] ),
    .A2(\w[50][19] ),
    .A3(\w[54][19] ),
    .S0(net502),
    .S1(net508),
    .X(_03002_));
 sky130_fd_sc_hd__mux4_2 _26250_ (.A0(\w[56][19] ),
    .A1(\w[60][19] ),
    .A2(\w[58][19] ),
    .A3(\w[62][19] ),
    .S0(net502),
    .S1(net508),
    .X(_03003_));
 sky130_fd_sc_hd__mux4_2 _26251_ (.A0(_03000_),
    .A1(_03001_),
    .A2(_03002_),
    .A3(_03003_),
    .S0(net497),
    .S1(net495),
    .X(_03004_));
 sky130_fd_sc_hd__mux2i_4 _26252_ (.A0(_02999_),
    .A1(_03004_),
    .S(net492),
    .Y(_03005_));
 sky130_fd_sc_hd__xnor2_1 _26253_ (.A(_02994_),
    .B(_03005_),
    .Y(_03006_));
 sky130_fd_sc_hd__xnor2_1 _26254_ (.A(_02976_),
    .B(_03006_),
    .Y(_11833_));
 sky130_fd_sc_hd__mux4_2 _26255_ (.A0(\w[0][1] ),
    .A1(\w[4][1] ),
    .A2(\w[2][1] ),
    .A3(\w[6][1] ),
    .S0(net381),
    .S1(net389),
    .X(_03007_));
 sky130_fd_sc_hd__mux4_2 _26256_ (.A0(\w[8][1] ),
    .A1(\w[12][1] ),
    .A2(\w[10][1] ),
    .A3(\w[14][1] ),
    .S0(net381),
    .S1(net389),
    .X(_03008_));
 sky130_fd_sc_hd__mux4_2 _26257_ (.A0(\w[16][1] ),
    .A1(\w[20][1] ),
    .A2(\w[18][1] ),
    .A3(\w[22][1] ),
    .S0(net381),
    .S1(net389),
    .X(_03009_));
 sky130_fd_sc_hd__mux4_2 _26258_ (.A0(\w[24][1] ),
    .A1(\w[28][1] ),
    .A2(\w[26][1] ),
    .A3(\w[30][1] ),
    .S0(net381),
    .S1(net389),
    .X(_03010_));
 sky130_fd_sc_hd__mux4_2 _26259_ (.A0(_03007_),
    .A1(_03008_),
    .A2(_03009_),
    .A3(_03010_),
    .S0(net378),
    .S1(net535),
    .X(_03011_));
 sky130_fd_sc_hd__mux4_2 _26260_ (.A0(\w[32][1] ),
    .A1(\w[36][1] ),
    .A2(\w[34][1] ),
    .A3(\w[38][1] ),
    .S0(net385),
    .S1(net392),
    .X(_03012_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_112 ();
 sky130_fd_sc_hd__mux4_2 _26262_ (.A0(\w[40][1] ),
    .A1(\w[44][1] ),
    .A2(\w[42][1] ),
    .A3(\w[46][1] ),
    .S0(net385),
    .S1(net392),
    .X(_03014_));
 sky130_fd_sc_hd__mux4_2 _26263_ (.A0(\w[48][1] ),
    .A1(\w[52][1] ),
    .A2(\w[50][1] ),
    .A3(\w[54][1] ),
    .S0(net385),
    .S1(net392),
    .X(_03015_));
 sky130_fd_sc_hd__mux4_2 _26264_ (.A0(\w[56][1] ),
    .A1(\w[60][1] ),
    .A2(\w[58][1] ),
    .A3(\w[62][1] ),
    .S0(net385),
    .S1(net392),
    .X(_03016_));
 sky130_fd_sc_hd__mux4_2 _26265_ (.A0(_03012_),
    .A1(_03014_),
    .A2(_03015_),
    .A3(_03016_),
    .S0(net378),
    .S1(net535),
    .X(_03017_));
 sky130_fd_sc_hd__mux2i_4 _26266_ (.A0(_03011_),
    .A1(_03017_),
    .S(net374),
    .Y(_11832_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 ();
 sky130_fd_sc_hd__mux4_2 _26275_ (.A0(\w[1][1] ),
    .A1(\w[5][1] ),
    .A2(\w[3][1] ),
    .A3(\w[7][1] ),
    .S0(net459),
    .S1(net470),
    .X(_03026_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 ();
 sky130_fd_sc_hd__mux4_2 _26280_ (.A0(\w[9][1] ),
    .A1(\w[13][1] ),
    .A2(\w[11][1] ),
    .A3(\w[15][1] ),
    .S0(net459),
    .S1(net544),
    .X(_03031_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_98 ();
 sky130_fd_sc_hd__mux4_2 _26283_ (.A0(\w[17][1] ),
    .A1(\w[21][1] ),
    .A2(\w[19][1] ),
    .A3(\w[23][1] ),
    .S0(net459),
    .S1(net470),
    .X(_03034_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_95 ();
 sky130_fd_sc_hd__mux4_2 _26287_ (.A0(\w[25][1] ),
    .A1(\w[29][1] ),
    .A2(\w[27][1] ),
    .A3(\w[31][1] ),
    .S0(net459),
    .S1(net470),
    .X(_03038_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_90 ();
 sky130_fd_sc_hd__mux4_2 _26293_ (.A0(_03026_),
    .A1(_03031_),
    .A2(_03034_),
    .A3(_03038_),
    .S0(net456),
    .S1(net454),
    .X(_03044_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_88 ();
 sky130_fd_sc_hd__mux4_2 _26296_ (.A0(\w[33][1] ),
    .A1(\w[37][1] ),
    .A2(\w[35][1] ),
    .A3(\w[39][1] ),
    .S0(net459),
    .S1(net470),
    .X(_03047_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_86 ();
 sky130_fd_sc_hd__mux4_2 _26299_ (.A0(\w[41][1] ),
    .A1(\w[45][1] ),
    .A2(\w[43][1] ),
    .A3(\w[47][1] ),
    .S0(net459),
    .S1(net470),
    .X(_03050_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_84 ();
 sky130_fd_sc_hd__mux4_2 _26302_ (.A0(\w[49][1] ),
    .A1(\w[53][1] ),
    .A2(\w[51][1] ),
    .A3(\w[55][1] ),
    .S0(net459),
    .S1(net470),
    .X(_03053_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_82 ();
 sky130_fd_sc_hd__mux4_2 _26305_ (.A0(\w[57][1] ),
    .A1(\w[61][1] ),
    .A2(\w[59][1] ),
    .A3(\w[63][1] ),
    .S0(net459),
    .S1(net470),
    .X(_03056_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_80 ();
 sky130_fd_sc_hd__mux4_2 _26308_ (.A0(_03047_),
    .A1(_03050_),
    .A2(_03053_),
    .A3(_03056_),
    .S0(net456),
    .S1(net454),
    .X(_03059_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_78 ();
 sky130_fd_sc_hd__mux2i_4 _26311_ (.A0(_03044_),
    .A1(_03059_),
    .S(net453),
    .Y(_11837_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_77 ();
 sky130_fd_sc_hd__mux4_2 _26313_ (.A0(\w[1][12] ),
    .A1(\w[5][12] ),
    .A2(\w[3][12] ),
    .A3(\w[7][12] ),
    .S0(net420),
    .S1(net427),
    .X(_03063_));
 sky130_fd_sc_hd__mux4_2 _26314_ (.A0(\w[9][12] ),
    .A1(\w[13][12] ),
    .A2(\w[11][12] ),
    .A3(\w[15][12] ),
    .S0(net420),
    .S1(net427),
    .X(_03064_));
 sky130_fd_sc_hd__mux4_2 _26315_ (.A0(\w[17][12] ),
    .A1(\w[21][12] ),
    .A2(\w[19][12] ),
    .A3(\w[23][12] ),
    .S0(net420),
    .S1(net427),
    .X(_03065_));
 sky130_fd_sc_hd__mux4_2 _26316_ (.A0(\w[25][12] ),
    .A1(\w[29][12] ),
    .A2(\w[27][12] ),
    .A3(\w[31][12] ),
    .S0(net420),
    .S1(net427),
    .X(_03066_));
 sky130_fd_sc_hd__mux4_2 _26317_ (.A0(_03063_),
    .A1(_03064_),
    .A2(_03065_),
    .A3(_03066_),
    .S0(net417),
    .S1(net415),
    .X(_03067_));
 sky130_fd_sc_hd__mux4_2 _26318_ (.A0(\w[33][12] ),
    .A1(\w[37][12] ),
    .A2(\w[35][12] ),
    .A3(\w[39][12] ),
    .S0(net421),
    .S1(net428),
    .X(_03068_));
 sky130_fd_sc_hd__mux4_2 _26319_ (.A0(\w[41][12] ),
    .A1(\w[45][12] ),
    .A2(\w[43][12] ),
    .A3(\w[47][12] ),
    .S0(net421),
    .S1(net428),
    .X(_03069_));
 sky130_fd_sc_hd__mux4_2 _26320_ (.A0(\w[49][12] ),
    .A1(\w[53][12] ),
    .A2(\w[51][12] ),
    .A3(\w[55][12] ),
    .S0(net421),
    .S1(net428),
    .X(_03070_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_76 ();
 sky130_fd_sc_hd__mux4_2 _26322_ (.A0(\w[57][12] ),
    .A1(\w[61][12] ),
    .A2(\w[59][12] ),
    .A3(\w[63][12] ),
    .S0(net421),
    .S1(net428),
    .X(_03072_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_75 ();
 sky130_fd_sc_hd__mux4_2 _26324_ (.A0(_03068_),
    .A1(_03069_),
    .A2(_03070_),
    .A3(_03072_),
    .S0(net418),
    .S1(net415),
    .X(_03074_));
 sky130_fd_sc_hd__mux2i_4 _26325_ (.A0(_03067_),
    .A1(_03074_),
    .S(net539),
    .Y(_03075_));
 sky130_fd_sc_hd__mux4_2 _26326_ (.A0(\w[1][21] ),
    .A1(\w[5][21] ),
    .A2(\w[3][21] ),
    .A3(\w[7][21] ),
    .S0(net420),
    .S1(net427),
    .X(_03076_));
 sky130_fd_sc_hd__mux4_2 _26327_ (.A0(\w[9][21] ),
    .A1(\w[13][21] ),
    .A2(\w[11][21] ),
    .A3(\w[15][21] ),
    .S0(net420),
    .S1(net427),
    .X(_03077_));
 sky130_fd_sc_hd__mux4_2 _26328_ (.A0(\w[17][21] ),
    .A1(\w[21][21] ),
    .A2(\w[19][21] ),
    .A3(\w[23][21] ),
    .S0(net420),
    .S1(net427),
    .X(_03078_));
 sky130_fd_sc_hd__mux4_2 _26329_ (.A0(\w[25][21] ),
    .A1(\w[29][21] ),
    .A2(\w[27][21] ),
    .A3(\w[31][21] ),
    .S0(net420),
    .S1(net427),
    .X(_03079_));
 sky130_fd_sc_hd__mux4_2 _26330_ (.A0(_03076_),
    .A1(_03077_),
    .A2(_03078_),
    .A3(_03079_),
    .S0(net418),
    .S1(net415),
    .X(_03080_));
 sky130_fd_sc_hd__mux4_2 _26331_ (.A0(\w[33][21] ),
    .A1(\w[37][21] ),
    .A2(\w[35][21] ),
    .A3(\w[39][21] ),
    .S0(net419),
    .S1(net426),
    .X(_03081_));
 sky130_fd_sc_hd__mux4_2 _26332_ (.A0(\w[41][21] ),
    .A1(\w[45][21] ),
    .A2(\w[43][21] ),
    .A3(\w[47][21] ),
    .S0(net419),
    .S1(net426),
    .X(_03082_));
 sky130_fd_sc_hd__mux4_2 _26333_ (.A0(\w[49][21] ),
    .A1(\w[53][21] ),
    .A2(\w[51][21] ),
    .A3(\w[55][21] ),
    .S0(net419),
    .S1(net426),
    .X(_03083_));
 sky130_fd_sc_hd__mux4_2 _26334_ (.A0(\w[57][21] ),
    .A1(\w[61][21] ),
    .A2(\w[59][21] ),
    .A3(\w[63][21] ),
    .S0(net419),
    .S1(net426),
    .X(_03084_));
 sky130_fd_sc_hd__mux4_2 _26335_ (.A0(_03081_),
    .A1(_03082_),
    .A2(_03083_),
    .A3(_03084_),
    .S0(net418),
    .S1(net415),
    .X(_03085_));
 sky130_fd_sc_hd__mux2i_4 _26336_ (.A0(_03080_),
    .A1(_03085_),
    .S(net539),
    .Y(_03086_));
 sky130_fd_sc_hd__xnor2_1 _26337_ (.A(_03075_),
    .B(_03086_),
    .Y(_03087_));
 sky130_fd_sc_hd__xnor2_1 _26338_ (.A(_02770_),
    .B(_03087_),
    .Y(_11842_));
 sky130_fd_sc_hd__mux4_2 _26339_ (.A0(\w[0][5] ),
    .A1(\w[4][5] ),
    .A2(\w[2][5] ),
    .A3(\w[6][5] ),
    .S0(\count15_2[2] ),
    .S1(net506),
    .X(_03088_));
 sky130_fd_sc_hd__mux4_2 _26340_ (.A0(\w[8][5] ),
    .A1(\w[12][5] ),
    .A2(\w[10][5] ),
    .A3(\w[14][5] ),
    .S0(\count15_2[2] ),
    .S1(net506),
    .X(_03089_));
 sky130_fd_sc_hd__mux4_2 _26341_ (.A0(\w[16][5] ),
    .A1(\w[20][5] ),
    .A2(\w[18][5] ),
    .A3(\w[22][5] ),
    .S0(\count15_2[2] ),
    .S1(net506),
    .X(_03090_));
 sky130_fd_sc_hd__mux4_2 _26342_ (.A0(\w[24][5] ),
    .A1(\w[28][5] ),
    .A2(\w[26][5] ),
    .A3(\w[30][5] ),
    .S0(\count15_2[2] ),
    .S1(net506),
    .X(_03091_));
 sky130_fd_sc_hd__mux4_2 _26343_ (.A0(_03088_),
    .A1(_03089_),
    .A2(_03090_),
    .A3(_03091_),
    .S0(net496),
    .S1(net547),
    .X(_03092_));
 sky130_fd_sc_hd__mux4_2 _26344_ (.A0(\w[32][5] ),
    .A1(\w[36][5] ),
    .A2(\w[34][5] ),
    .A3(\w[38][5] ),
    .S0(net499),
    .S1(net506),
    .X(_03093_));
 sky130_fd_sc_hd__mux4_2 _26345_ (.A0(\w[40][5] ),
    .A1(\w[44][5] ),
    .A2(\w[42][5] ),
    .A3(\w[46][5] ),
    .S0(net499),
    .S1(net506),
    .X(_03094_));
 sky130_fd_sc_hd__mux4_2 _26346_ (.A0(\w[48][5] ),
    .A1(\w[52][5] ),
    .A2(\w[50][5] ),
    .A3(\w[54][5] ),
    .S0(net499),
    .S1(net506),
    .X(_03095_));
 sky130_fd_sc_hd__mux4_2 _26347_ (.A0(\w[56][5] ),
    .A1(\w[60][5] ),
    .A2(\w[58][5] ),
    .A3(\w[62][5] ),
    .S0(net499),
    .S1(net506),
    .X(_03096_));
 sky130_fd_sc_hd__mux4_2 _26348_ (.A0(_03093_),
    .A1(_03094_),
    .A2(_03095_),
    .A3(_03096_),
    .S0(net496),
    .S1(net547),
    .X(_03097_));
 sky130_fd_sc_hd__mux2i_4 _26349_ (.A0(_03092_),
    .A1(_03097_),
    .S(net493),
    .Y(_03098_));
 sky130_fd_sc_hd__mux4_2 _26350_ (.A0(\w[0][20] ),
    .A1(\w[4][20] ),
    .A2(\w[2][20] ),
    .A3(\w[6][20] ),
    .S0(net502),
    .S1(net508),
    .X(_03099_));
 sky130_fd_sc_hd__mux4_2 _26351_ (.A0(\w[8][20] ),
    .A1(\w[12][20] ),
    .A2(\w[10][20] ),
    .A3(\w[14][20] ),
    .S0(net502),
    .S1(net508),
    .X(_03100_));
 sky130_fd_sc_hd__mux4_2 _26352_ (.A0(\w[16][20] ),
    .A1(\w[20][20] ),
    .A2(\w[18][20] ),
    .A3(\w[22][20] ),
    .S0(net502),
    .S1(net508),
    .X(_03101_));
 sky130_fd_sc_hd__mux4_2 _26353_ (.A0(\w[24][20] ),
    .A1(\w[28][20] ),
    .A2(\w[26][20] ),
    .A3(\w[30][20] ),
    .S0(net502),
    .S1(net508),
    .X(_03102_));
 sky130_fd_sc_hd__mux4_2 _26354_ (.A0(_03099_),
    .A1(_03100_),
    .A2(_03101_),
    .A3(_03102_),
    .S0(net497),
    .S1(net495),
    .X(_03103_));
 sky130_fd_sc_hd__mux4_2 _26355_ (.A0(\w[32][20] ),
    .A1(\w[36][20] ),
    .A2(\w[34][20] ),
    .A3(\w[38][20] ),
    .S0(net504),
    .S1(net510),
    .X(_03104_));
 sky130_fd_sc_hd__mux4_2 _26356_ (.A0(\w[40][20] ),
    .A1(\w[44][20] ),
    .A2(\w[42][20] ),
    .A3(\w[46][20] ),
    .S0(net504),
    .S1(net510),
    .X(_03105_));
 sky130_fd_sc_hd__mux4_2 _26357_ (.A0(\w[48][20] ),
    .A1(\w[52][20] ),
    .A2(\w[50][20] ),
    .A3(\w[54][20] ),
    .S0(net504),
    .S1(net510),
    .X(_03106_));
 sky130_fd_sc_hd__mux4_2 _26358_ (.A0(\w[56][20] ),
    .A1(\w[60][20] ),
    .A2(\w[58][20] ),
    .A3(\w[62][20] ),
    .S0(net504),
    .S1(net510),
    .X(_03107_));
 sky130_fd_sc_hd__mux4_2 _26359_ (.A0(_03104_),
    .A1(_03105_),
    .A2(_03106_),
    .A3(_03107_),
    .S0(net497),
    .S1(net495),
    .X(_03108_));
 sky130_fd_sc_hd__mux2i_4 _26360_ (.A0(_03103_),
    .A1(_03108_),
    .S(net492),
    .Y(_03109_));
 sky130_fd_sc_hd__mux4_2 _26361_ (.A0(\w[0][9] ),
    .A1(\w[4][9] ),
    .A2(\w[2][9] ),
    .A3(\w[6][9] ),
    .S0(net500),
    .S1(net507),
    .X(_03110_));
 sky130_fd_sc_hd__mux4_2 _26362_ (.A0(\w[8][9] ),
    .A1(\w[12][9] ),
    .A2(\w[10][9] ),
    .A3(\w[14][9] ),
    .S0(net500),
    .S1(net507),
    .X(_03111_));
 sky130_fd_sc_hd__mux4_2 _26363_ (.A0(\w[16][9] ),
    .A1(\w[20][9] ),
    .A2(\w[18][9] ),
    .A3(\w[22][9] ),
    .S0(net500),
    .S1(net507),
    .X(_03112_));
 sky130_fd_sc_hd__mux4_2 _26364_ (.A0(\w[24][9] ),
    .A1(\w[28][9] ),
    .A2(\w[26][9] ),
    .A3(\w[30][9] ),
    .S0(net500),
    .S1(net507),
    .X(_03113_));
 sky130_fd_sc_hd__mux4_2 _26365_ (.A0(_03110_),
    .A1(_03111_),
    .A2(_03112_),
    .A3(_03113_),
    .S0(net497),
    .S1(net495),
    .X(_03114_));
 sky130_fd_sc_hd__mux4_2 _26366_ (.A0(\w[32][9] ),
    .A1(\w[36][9] ),
    .A2(\w[34][9] ),
    .A3(\w[38][9] ),
    .S0(net502),
    .S1(net508),
    .X(_03115_));
 sky130_fd_sc_hd__mux4_2 _26367_ (.A0(\w[40][9] ),
    .A1(\w[44][9] ),
    .A2(\w[42][9] ),
    .A3(\w[46][9] ),
    .S0(net502),
    .S1(net508),
    .X(_03116_));
 sky130_fd_sc_hd__mux4_2 _26368_ (.A0(\w[48][9] ),
    .A1(\w[52][9] ),
    .A2(\w[50][9] ),
    .A3(\w[54][9] ),
    .S0(net502),
    .S1(net508),
    .X(_03117_));
 sky130_fd_sc_hd__mux4_2 _26369_ (.A0(\w[56][9] ),
    .A1(\w[60][9] ),
    .A2(\w[58][9] ),
    .A3(\w[62][9] ),
    .S0(net502),
    .S1(net508),
    .X(_03118_));
 sky130_fd_sc_hd__mux4_2 _26370_ (.A0(_03115_),
    .A1(_03116_),
    .A2(_03117_),
    .A3(_03118_),
    .S0(net548),
    .S1(net494),
    .X(_03119_));
 sky130_fd_sc_hd__mux2i_4 _26371_ (.A0(_03114_),
    .A1(_03119_),
    .S(net492),
    .Y(_03120_));
 sky130_fd_sc_hd__xnor2_1 _26372_ (.A(_03109_),
    .B(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__xnor2_1 _26373_ (.A(_03098_),
    .B(_03121_),
    .Y(_11841_));
 sky130_fd_sc_hd__mux4_2 _26374_ (.A0(\w[0][2] ),
    .A1(\w[4][2] ),
    .A2(\w[2][2] ),
    .A3(\w[6][2] ),
    .S0(net380),
    .S1(net388),
    .X(_03122_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_74 ();
 sky130_fd_sc_hd__mux4_2 _26376_ (.A0(\w[8][2] ),
    .A1(\w[12][2] ),
    .A2(\w[10][2] ),
    .A3(\w[14][2] ),
    .S0(net380),
    .S1(net388),
    .X(_03124_));
 sky130_fd_sc_hd__mux4_2 _26377_ (.A0(\w[16][2] ),
    .A1(\w[20][2] ),
    .A2(\w[18][2] ),
    .A3(\w[22][2] ),
    .S0(net380),
    .S1(net388),
    .X(_03125_));
 sky130_fd_sc_hd__mux4_2 _26378_ (.A0(\w[24][2] ),
    .A1(\w[28][2] ),
    .A2(\w[26][2] ),
    .A3(\w[30][2] ),
    .S0(net380),
    .S1(net388),
    .X(_03126_));
 sky130_fd_sc_hd__mux4_2 _26379_ (.A0(_03122_),
    .A1(_03124_),
    .A2(_03125_),
    .A3(_03126_),
    .S0(net379),
    .S1(net376),
    .X(_03127_));
 sky130_fd_sc_hd__mux4_2 _26380_ (.A0(\w[32][2] ),
    .A1(\w[36][2] ),
    .A2(\w[34][2] ),
    .A3(\w[38][2] ),
    .S0(net386),
    .S1(net393),
    .X(_03128_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_73 ();
 sky130_fd_sc_hd__mux4_2 _26382_ (.A0(\w[40][2] ),
    .A1(\w[44][2] ),
    .A2(\w[42][2] ),
    .A3(\w[46][2] ),
    .S0(net386),
    .S1(net393),
    .X(_03130_));
 sky130_fd_sc_hd__mux4_2 _26383_ (.A0(\w[48][2] ),
    .A1(\w[52][2] ),
    .A2(\w[50][2] ),
    .A3(\w[54][2] ),
    .S0(net386),
    .S1(net393),
    .X(_03131_));
 sky130_fd_sc_hd__mux4_2 _26384_ (.A0(\w[56][2] ),
    .A1(\w[60][2] ),
    .A2(\w[58][2] ),
    .A3(\w[62][2] ),
    .S0(net386),
    .S1(net393),
    .X(_03132_));
 sky130_fd_sc_hd__mux4_2 _26385_ (.A0(_03128_),
    .A1(_03130_),
    .A2(_03131_),
    .A3(_03132_),
    .S0(net379),
    .S1(net376),
    .X(_03133_));
 sky130_fd_sc_hd__mux2i_4 _26386_ (.A0(_03127_),
    .A1(_03133_),
    .S(net373),
    .Y(_11840_));
 sky130_fd_sc_hd__mux4_2 _26387_ (.A0(\w[1][2] ),
    .A1(\w[5][2] ),
    .A2(\w[3][2] ),
    .A3(\w[7][2] ),
    .S0(net460),
    .S1(net470),
    .X(_03134_));
 sky130_fd_sc_hd__mux4_2 _26388_ (.A0(\w[9][2] ),
    .A1(\w[13][2] ),
    .A2(\w[11][2] ),
    .A3(\w[15][2] ),
    .S0(net460),
    .S1(net470),
    .X(_03135_));
 sky130_fd_sc_hd__mux4_2 _26389_ (.A0(\w[17][2] ),
    .A1(\w[21][2] ),
    .A2(\w[19][2] ),
    .A3(\w[23][2] ),
    .S0(net460),
    .S1(net470),
    .X(_03136_));
 sky130_fd_sc_hd__mux4_2 _26390_ (.A0(\w[25][2] ),
    .A1(\w[29][2] ),
    .A2(\w[27][2] ),
    .A3(\w[31][2] ),
    .S0(net460),
    .S1(net470),
    .X(_03137_));
 sky130_fd_sc_hd__mux4_2 _26391_ (.A0(_03134_),
    .A1(_03135_),
    .A2(_03136_),
    .A3(_03137_),
    .S0(net456),
    .S1(net454),
    .X(_03138_));
 sky130_fd_sc_hd__mux4_2 _26392_ (.A0(\w[33][2] ),
    .A1(\w[37][2] ),
    .A2(\w[35][2] ),
    .A3(\w[39][2] ),
    .S0(net460),
    .S1(net468),
    .X(_03139_));
 sky130_fd_sc_hd__mux4_2 _26393_ (.A0(\w[41][2] ),
    .A1(\w[45][2] ),
    .A2(\w[43][2] ),
    .A3(\w[47][2] ),
    .S0(net460),
    .S1(net468),
    .X(_03140_));
 sky130_fd_sc_hd__mux4_2 _26394_ (.A0(\w[49][2] ),
    .A1(\w[53][2] ),
    .A2(\w[51][2] ),
    .A3(\w[55][2] ),
    .S0(net460),
    .S1(net468),
    .X(_03141_));
 sky130_fd_sc_hd__mux4_2 _26395_ (.A0(\w[57][2] ),
    .A1(\w[61][2] ),
    .A2(\w[59][2] ),
    .A3(\w[63][2] ),
    .S0(net460),
    .S1(net468),
    .X(_03142_));
 sky130_fd_sc_hd__mux4_2 _26396_ (.A0(_03139_),
    .A1(_03140_),
    .A2(_03141_),
    .A3(_03142_),
    .S0(net456),
    .S1(net454),
    .X(_03143_));
 sky130_fd_sc_hd__mux2i_4 _26397_ (.A0(_03138_),
    .A1(_03143_),
    .S(net453),
    .Y(_11845_));
 sky130_fd_sc_hd__mux4_2 _26398_ (.A0(\w[1][13] ),
    .A1(\w[5][13] ),
    .A2(\w[3][13] ),
    .A3(\w[7][13] ),
    .S0(net419),
    .S1(net426),
    .X(_03144_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_71 ();
 sky130_fd_sc_hd__mux4_2 _26401_ (.A0(\w[9][13] ),
    .A1(\w[13][13] ),
    .A2(\w[11][13] ),
    .A3(\w[15][13] ),
    .S0(net419),
    .S1(net426),
    .X(_03147_));
 sky130_fd_sc_hd__mux4_2 _26402_ (.A0(\w[17][13] ),
    .A1(\w[21][13] ),
    .A2(\w[19][13] ),
    .A3(\w[23][13] ),
    .S0(net419),
    .S1(net426),
    .X(_03148_));
 sky130_fd_sc_hd__mux4_2 _26403_ (.A0(\w[25][13] ),
    .A1(\w[29][13] ),
    .A2(\w[27][13] ),
    .A3(\w[31][13] ),
    .S0(net419),
    .S1(net426),
    .X(_03149_));
 sky130_fd_sc_hd__mux4_2 _26404_ (.A0(_03144_),
    .A1(_03147_),
    .A2(_03148_),
    .A3(_03149_),
    .S0(net418),
    .S1(net415),
    .X(_03150_));
 sky130_fd_sc_hd__mux4_2 _26405_ (.A0(\w[33][13] ),
    .A1(\w[37][13] ),
    .A2(\w[35][13] ),
    .A3(\w[39][13] ),
    .S0(net425),
    .S1(net430),
    .X(_03151_));
 sky130_fd_sc_hd__mux4_2 _26406_ (.A0(\w[41][13] ),
    .A1(\w[45][13] ),
    .A2(\w[43][13] ),
    .A3(\w[47][13] ),
    .S0(net425),
    .S1(net430),
    .X(_03152_));
 sky130_fd_sc_hd__mux4_2 _26407_ (.A0(\w[49][13] ),
    .A1(\w[53][13] ),
    .A2(\w[51][13] ),
    .A3(\w[55][13] ),
    .S0(net425),
    .S1(net430),
    .X(_03153_));
 sky130_fd_sc_hd__mux4_2 _26408_ (.A0(\w[57][13] ),
    .A1(\w[61][13] ),
    .A2(\w[59][13] ),
    .A3(\w[63][13] ),
    .S0(net425),
    .S1(net430),
    .X(_03154_));
 sky130_fd_sc_hd__mux4_2 _26409_ (.A0(_03151_),
    .A1(_03152_),
    .A2(_03153_),
    .A3(_03154_),
    .S0(net418),
    .S1(net415),
    .X(_03155_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_70 ();
 sky130_fd_sc_hd__mux2i_4 _26411_ (.A0(_03150_),
    .A1(_03155_),
    .S(net539),
    .Y(_03157_));
 sky130_fd_sc_hd__mux4_2 _26412_ (.A0(\w[1][22] ),
    .A1(\w[5][22] ),
    .A2(\w[3][22] ),
    .A3(\w[7][22] ),
    .S0(net420),
    .S1(net427),
    .X(_03158_));
 sky130_fd_sc_hd__mux4_2 _26413_ (.A0(\w[9][22] ),
    .A1(\w[13][22] ),
    .A2(\w[11][22] ),
    .A3(\w[15][22] ),
    .S0(net420),
    .S1(net427),
    .X(_03159_));
 sky130_fd_sc_hd__mux4_2 _26414_ (.A0(\w[17][22] ),
    .A1(\w[21][22] ),
    .A2(\w[19][22] ),
    .A3(\w[23][22] ),
    .S0(net420),
    .S1(net427),
    .X(_03160_));
 sky130_fd_sc_hd__mux4_2 _26415_ (.A0(\w[25][22] ),
    .A1(\w[29][22] ),
    .A2(\w[27][22] ),
    .A3(\w[31][22] ),
    .S0(net420),
    .S1(net427),
    .X(_03161_));
 sky130_fd_sc_hd__mux4_2 _26416_ (.A0(_03158_),
    .A1(_03159_),
    .A2(_03160_),
    .A3(_03161_),
    .S0(net416),
    .S1(net415),
    .X(_03162_));
 sky130_fd_sc_hd__mux4_2 _26417_ (.A0(\w[33][22] ),
    .A1(\w[37][22] ),
    .A2(\w[35][22] ),
    .A3(\w[39][22] ),
    .S0(net420),
    .S1(net427),
    .X(_03163_));
 sky130_fd_sc_hd__mux4_2 _26418_ (.A0(\w[41][22] ),
    .A1(\w[45][22] ),
    .A2(\w[43][22] ),
    .A3(\w[47][22] ),
    .S0(net420),
    .S1(net427),
    .X(_03164_));
 sky130_fd_sc_hd__mux4_2 _26419_ (.A0(\w[49][22] ),
    .A1(\w[53][22] ),
    .A2(\w[51][22] ),
    .A3(\w[55][22] ),
    .S0(net420),
    .S1(net427),
    .X(_03165_));
 sky130_fd_sc_hd__mux4_2 _26420_ (.A0(\w[57][22] ),
    .A1(\w[61][22] ),
    .A2(\w[59][22] ),
    .A3(\w[63][22] ),
    .S0(net420),
    .S1(net427),
    .X(_03166_));
 sky130_fd_sc_hd__mux4_2 _26421_ (.A0(_03163_),
    .A1(_03164_),
    .A2(_03165_),
    .A3(_03166_),
    .S0(net417),
    .S1(net415),
    .X(_03167_));
 sky130_fd_sc_hd__mux2i_4 _26422_ (.A0(_03162_),
    .A1(_03167_),
    .S(net413),
    .Y(_03168_));
 sky130_fd_sc_hd__xnor2_1 _26423_ (.A(_03157_),
    .B(_03168_),
    .Y(_03169_));
 sky130_fd_sc_hd__xnor2_1 _26424_ (.A(_02953_),
    .B(_03169_),
    .Y(_11853_));
 sky130_fd_sc_hd__mux4_2 _26425_ (.A0(\w[0][21] ),
    .A1(\w[4][21] ),
    .A2(\w[2][21] ),
    .A3(\w[6][21] ),
    .S0(net501),
    .S1(net507),
    .X(_03170_));
 sky130_fd_sc_hd__mux4_2 _26426_ (.A0(\w[8][21] ),
    .A1(\w[12][21] ),
    .A2(\w[10][21] ),
    .A3(\w[14][21] ),
    .S0(net501),
    .S1(net507),
    .X(_03171_));
 sky130_fd_sc_hd__mux4_2 _26427_ (.A0(\w[16][21] ),
    .A1(\w[20][21] ),
    .A2(\w[18][21] ),
    .A3(\w[22][21] ),
    .S0(net501),
    .S1(net507),
    .X(_03172_));
 sky130_fd_sc_hd__mux4_2 _26428_ (.A0(\w[24][21] ),
    .A1(\w[28][21] ),
    .A2(\w[26][21] ),
    .A3(\w[30][21] ),
    .S0(net501),
    .S1(net507),
    .X(_03173_));
 sky130_fd_sc_hd__mux4_2 _26429_ (.A0(_03170_),
    .A1(_03171_),
    .A2(_03172_),
    .A3(_03173_),
    .S0(net548),
    .S1(net494),
    .X(_03174_));
 sky130_fd_sc_hd__mux4_2 _26430_ (.A0(\w[32][21] ),
    .A1(\w[36][21] ),
    .A2(\w[34][21] ),
    .A3(\w[38][21] ),
    .S0(net504),
    .S1(net510),
    .X(_03175_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_69 ();
 sky130_fd_sc_hd__mux4_2 _26432_ (.A0(\w[40][21] ),
    .A1(\w[44][21] ),
    .A2(\w[42][21] ),
    .A3(\w[46][21] ),
    .S0(net504),
    .S1(net510),
    .X(_03177_));
 sky130_fd_sc_hd__mux4_2 _26433_ (.A0(\w[48][21] ),
    .A1(\w[52][21] ),
    .A2(\w[50][21] ),
    .A3(\w[54][21] ),
    .S0(net504),
    .S1(net510),
    .X(_03178_));
 sky130_fd_sc_hd__mux4_2 _26434_ (.A0(\w[56][21] ),
    .A1(\w[60][21] ),
    .A2(\w[58][21] ),
    .A3(\w[62][21] ),
    .S0(net504),
    .S1(net510),
    .X(_03179_));
 sky130_fd_sc_hd__mux4_2 _26435_ (.A0(_03175_),
    .A1(_03177_),
    .A2(_03178_),
    .A3(_03179_),
    .S0(net548),
    .S1(net494),
    .X(_03180_));
 sky130_fd_sc_hd__mux2i_4 _26436_ (.A0(_03174_),
    .A1(_03180_),
    .S(net492),
    .Y(_03181_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_67 ();
 sky130_fd_sc_hd__mux4_2 _26439_ (.A0(\w[0][6] ),
    .A1(\w[4][6] ),
    .A2(\w[2][6] ),
    .A3(\w[6][6] ),
    .S0(\count15_2[2] ),
    .S1(net506),
    .X(_03184_));
 sky130_fd_sc_hd__mux4_2 _26440_ (.A0(\w[8][6] ),
    .A1(\w[12][6] ),
    .A2(\w[10][6] ),
    .A3(\w[14][6] ),
    .S0(\count15_2[2] ),
    .S1(net506),
    .X(_03185_));
 sky130_fd_sc_hd__mux4_2 _26441_ (.A0(\w[16][6] ),
    .A1(\w[20][6] ),
    .A2(\w[18][6] ),
    .A3(\w[22][6] ),
    .S0(\count15_2[2] ),
    .S1(net506),
    .X(_03186_));
 sky130_fd_sc_hd__mux4_2 _26442_ (.A0(\w[24][6] ),
    .A1(\w[28][6] ),
    .A2(\w[26][6] ),
    .A3(\w[30][6] ),
    .S0(net499),
    .S1(net506),
    .X(_03187_));
 sky130_fd_sc_hd__mux4_2 _26443_ (.A0(_03184_),
    .A1(_03185_),
    .A2(_03186_),
    .A3(_03187_),
    .S0(\count15_2[3] ),
    .S1(net547),
    .X(_03188_));
 sky130_fd_sc_hd__mux4_2 _26444_ (.A0(\w[32][6] ),
    .A1(\w[36][6] ),
    .A2(\w[34][6] ),
    .A3(\w[38][6] ),
    .S0(net505),
    .S1(\count15_2[1] ),
    .X(_03189_));
 sky130_fd_sc_hd__mux4_2 _26445_ (.A0(\w[40][6] ),
    .A1(\w[44][6] ),
    .A2(\w[42][6] ),
    .A3(\w[46][6] ),
    .S0(net505),
    .S1(\count15_2[1] ),
    .X(_03190_));
 sky130_fd_sc_hd__mux4_2 _26446_ (.A0(\w[48][6] ),
    .A1(\w[52][6] ),
    .A2(\w[50][6] ),
    .A3(\w[54][6] ),
    .S0(net505),
    .S1(\count15_2[1] ),
    .X(_03191_));
 sky130_fd_sc_hd__mux4_2 _26447_ (.A0(\w[56][6] ),
    .A1(\w[60][6] ),
    .A2(\w[58][6] ),
    .A3(\w[62][6] ),
    .S0(net505),
    .S1(\count15_2[1] ),
    .X(_03192_));
 sky130_fd_sc_hd__mux4_2 _26448_ (.A0(_03189_),
    .A1(_03190_),
    .A2(_03191_),
    .A3(_03192_),
    .S0(net497),
    .S1(\count15_2[4] ),
    .X(_03193_));
 sky130_fd_sc_hd__mux2i_4 _26449_ (.A0(_03188_),
    .A1(_03193_),
    .S(net493),
    .Y(_03194_));
 sky130_fd_sc_hd__mux4_2 _26450_ (.A0(\w[0][10] ),
    .A1(\w[4][10] ),
    .A2(\w[2][10] ),
    .A3(\w[6][10] ),
    .S0(net500),
    .S1(net507),
    .X(_03195_));
 sky130_fd_sc_hd__mux4_2 _26451_ (.A0(\w[8][10] ),
    .A1(\w[12][10] ),
    .A2(\w[10][10] ),
    .A3(\w[14][10] ),
    .S0(net500),
    .S1(net507),
    .X(_03196_));
 sky130_fd_sc_hd__mux4_2 _26452_ (.A0(\w[16][10] ),
    .A1(\w[20][10] ),
    .A2(\w[18][10] ),
    .A3(\w[22][10] ),
    .S0(net500),
    .S1(net507),
    .X(_03197_));
 sky130_fd_sc_hd__mux4_2 _26453_ (.A0(\w[24][10] ),
    .A1(\w[28][10] ),
    .A2(\w[26][10] ),
    .A3(\w[30][10] ),
    .S0(net500),
    .S1(net507),
    .X(_03198_));
 sky130_fd_sc_hd__mux4_2 _26454_ (.A0(_03195_),
    .A1(_03196_),
    .A2(_03197_),
    .A3(_03198_),
    .S0(net497),
    .S1(net495),
    .X(_03199_));
 sky130_fd_sc_hd__mux4_2 _26455_ (.A0(\w[32][10] ),
    .A1(\w[36][10] ),
    .A2(\w[34][10] ),
    .A3(\w[38][10] ),
    .S0(net502),
    .S1(net508),
    .X(_03200_));
 sky130_fd_sc_hd__mux4_2 _26456_ (.A0(\w[40][10] ),
    .A1(\w[44][10] ),
    .A2(\w[42][10] ),
    .A3(\w[46][10] ),
    .S0(net502),
    .S1(net508),
    .X(_03201_));
 sky130_fd_sc_hd__mux4_2 _26457_ (.A0(\w[48][10] ),
    .A1(\w[52][10] ),
    .A2(\w[50][10] ),
    .A3(\w[54][10] ),
    .S0(net502),
    .S1(net508),
    .X(_03202_));
 sky130_fd_sc_hd__mux4_2 _26458_ (.A0(\w[56][10] ),
    .A1(\w[60][10] ),
    .A2(\w[58][10] ),
    .A3(\w[62][10] ),
    .S0(net502),
    .S1(net508),
    .X(_03203_));
 sky130_fd_sc_hd__mux4_2 _26459_ (.A0(_03200_),
    .A1(_03201_),
    .A2(_03202_),
    .A3(_03203_),
    .S0(net497),
    .S1(net495),
    .X(_03204_));
 sky130_fd_sc_hd__mux2i_4 _26460_ (.A0(_03199_),
    .A1(_03204_),
    .S(net492),
    .Y(_03205_));
 sky130_fd_sc_hd__xnor2_1 _26461_ (.A(_03194_),
    .B(_03205_),
    .Y(_03206_));
 sky130_fd_sc_hd__xnor2_1 _26462_ (.A(_03181_),
    .B(_03206_),
    .Y(_11852_));
 sky130_fd_sc_hd__mux4_2 _26463_ (.A0(\w[0][3] ),
    .A1(\w[4][3] ),
    .A2(\w[2][3] ),
    .A3(\w[6][3] ),
    .S0(net387),
    .S1(\count7_2[1] ),
    .X(_03207_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_66 ();
 sky130_fd_sc_hd__mux4_2 _26465_ (.A0(\w[8][3] ),
    .A1(\w[12][3] ),
    .A2(\w[10][3] ),
    .A3(\w[14][3] ),
    .S0(net387),
    .S1(\count7_2[1] ),
    .X(_03209_));
 sky130_fd_sc_hd__mux4_2 _26466_ (.A0(\w[16][3] ),
    .A1(\w[20][3] ),
    .A2(\w[18][3] ),
    .A3(\w[22][3] ),
    .S0(net387),
    .S1(\count7_2[1] ),
    .X(_03210_));
 sky130_fd_sc_hd__mux4_2 _26467_ (.A0(\w[24][3] ),
    .A1(\w[28][3] ),
    .A2(\w[26][3] ),
    .A3(\w[30][3] ),
    .S0(net387),
    .S1(\count7_2[1] ),
    .X(_03211_));
 sky130_fd_sc_hd__mux4_2 _26468_ (.A0(_03207_),
    .A1(_03209_),
    .A2(_03210_),
    .A3(_03211_),
    .S0(\count7_2[3] ),
    .S1(net376),
    .X(_03212_));
 sky130_fd_sc_hd__mux4_2 _26469_ (.A0(\w[32][3] ),
    .A1(\w[36][3] ),
    .A2(\w[34][3] ),
    .A3(\w[38][3] ),
    .S0(net387),
    .S1(\count7_2[1] ),
    .X(_03213_));
 sky130_fd_sc_hd__mux4_2 _26470_ (.A0(\w[40][3] ),
    .A1(\w[44][3] ),
    .A2(\w[42][3] ),
    .A3(\w[46][3] ),
    .S0(net387),
    .S1(\count7_2[1] ),
    .X(_03214_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_65 ();
 sky130_fd_sc_hd__mux4_2 _26472_ (.A0(\w[48][3] ),
    .A1(\w[52][3] ),
    .A2(\w[50][3] ),
    .A3(\w[54][3] ),
    .S0(net387),
    .S1(\count7_2[1] ),
    .X(_03216_));
 sky130_fd_sc_hd__mux4_2 _26473_ (.A0(\w[56][3] ),
    .A1(\w[60][3] ),
    .A2(\w[58][3] ),
    .A3(\w[62][3] ),
    .S0(net387),
    .S1(net393),
    .X(_03217_));
 sky130_fd_sc_hd__mux4_2 _26474_ (.A0(_03213_),
    .A1(_03214_),
    .A2(_03216_),
    .A3(_03217_),
    .S0(\count7_2[3] ),
    .S1(net376),
    .X(_03218_));
 sky130_fd_sc_hd__mux2i_4 _26475_ (.A0(_03212_),
    .A1(_03218_),
    .S(\count7_2[5] ),
    .Y(_11851_));
 sky130_fd_sc_hd__mux4_2 _26476_ (.A0(\w[1][3] ),
    .A1(\w[5][3] ),
    .A2(\w[3][3] ),
    .A3(\w[7][3] ),
    .S0(net461),
    .S1(net544),
    .X(_03219_));
 sky130_fd_sc_hd__mux4_2 _26477_ (.A0(\w[9][3] ),
    .A1(\w[13][3] ),
    .A2(\w[11][3] ),
    .A3(\w[15][3] ),
    .S0(net461),
    .S1(net544),
    .X(_03220_));
 sky130_fd_sc_hd__mux4_2 _26478_ (.A0(\w[17][3] ),
    .A1(\w[21][3] ),
    .A2(\w[19][3] ),
    .A3(\w[23][3] ),
    .S0(net461),
    .S1(net544),
    .X(_03221_));
 sky130_fd_sc_hd__mux4_2 _26479_ (.A0(\w[25][3] ),
    .A1(\w[29][3] ),
    .A2(\w[27][3] ),
    .A3(\w[31][3] ),
    .S0(net461),
    .S1(net544),
    .X(_03222_));
 sky130_fd_sc_hd__mux4_2 _26480_ (.A0(_03219_),
    .A1(_03220_),
    .A2(_03221_),
    .A3(_03222_),
    .S0(net456),
    .S1(net454),
    .X(_03223_));
 sky130_fd_sc_hd__mux4_2 _26481_ (.A0(\w[33][3] ),
    .A1(\w[37][3] ),
    .A2(\w[35][3] ),
    .A3(\w[39][3] ),
    .S0(net461),
    .S1(net544),
    .X(_03224_));
 sky130_fd_sc_hd__mux4_2 _26482_ (.A0(\w[41][3] ),
    .A1(\w[45][3] ),
    .A2(\w[43][3] ),
    .A3(\w[47][3] ),
    .S0(net461),
    .S1(net544),
    .X(_03225_));
 sky130_fd_sc_hd__mux4_2 _26483_ (.A0(\w[49][3] ),
    .A1(\w[53][3] ),
    .A2(\w[51][3] ),
    .A3(\w[55][3] ),
    .S0(net461),
    .S1(net544),
    .X(_03226_));
 sky130_fd_sc_hd__mux4_2 _26484_ (.A0(\w[57][3] ),
    .A1(\w[61][3] ),
    .A2(\w[59][3] ),
    .A3(\w[63][3] ),
    .S0(net461),
    .S1(net544),
    .X(_03227_));
 sky130_fd_sc_hd__mux4_2 _26485_ (.A0(_03224_),
    .A1(_03225_),
    .A2(_03226_),
    .A3(_03227_),
    .S0(net457),
    .S1(net543),
    .X(_03228_));
 sky130_fd_sc_hd__mux2i_4 _26486_ (.A0(_03223_),
    .A1(_03228_),
    .S(net453),
    .Y(_11856_));
 sky130_fd_sc_hd__mux4_2 _26487_ (.A0(\w[1][14] ),
    .A1(\w[5][14] ),
    .A2(\w[3][14] ),
    .A3(\w[7][14] ),
    .S0(net423),
    .S1(net427),
    .X(_03229_));
 sky130_fd_sc_hd__mux4_2 _26488_ (.A0(\w[9][14] ),
    .A1(\w[13][14] ),
    .A2(\w[11][14] ),
    .A3(\w[15][14] ),
    .S0(net423),
    .S1(net427),
    .X(_03230_));
 sky130_fd_sc_hd__mux4_2 _26489_ (.A0(\w[17][14] ),
    .A1(\w[21][14] ),
    .A2(\w[19][14] ),
    .A3(\w[23][14] ),
    .S0(net423),
    .S1(net427),
    .X(_03231_));
 sky130_fd_sc_hd__mux4_2 _26490_ (.A0(\w[25][14] ),
    .A1(\w[29][14] ),
    .A2(\w[27][14] ),
    .A3(\w[31][14] ),
    .S0(net423),
    .S1(net427),
    .X(_03232_));
 sky130_fd_sc_hd__mux4_2 _26491_ (.A0(_03229_),
    .A1(_03230_),
    .A2(_03231_),
    .A3(_03232_),
    .S0(net416),
    .S1(net414),
    .X(_03233_));
 sky130_fd_sc_hd__mux4_2 _26492_ (.A0(\w[33][14] ),
    .A1(\w[37][14] ),
    .A2(\w[35][14] ),
    .A3(\w[39][14] ),
    .S0(net420),
    .S1(net427),
    .X(_03234_));
 sky130_fd_sc_hd__mux4_2 _26493_ (.A0(\w[41][14] ),
    .A1(\w[45][14] ),
    .A2(\w[43][14] ),
    .A3(\w[47][14] ),
    .S0(net420),
    .S1(net427),
    .X(_03235_));
 sky130_fd_sc_hd__mux4_2 _26494_ (.A0(\w[49][14] ),
    .A1(\w[53][14] ),
    .A2(\w[51][14] ),
    .A3(\w[55][14] ),
    .S0(net420),
    .S1(net427),
    .X(_03236_));
 sky130_fd_sc_hd__mux4_2 _26495_ (.A0(\w[57][14] ),
    .A1(\w[61][14] ),
    .A2(\w[59][14] ),
    .A3(\w[63][14] ),
    .S0(net420),
    .S1(net427),
    .X(_03237_));
 sky130_fd_sc_hd__mux4_2 _26496_ (.A0(_03234_),
    .A1(_03235_),
    .A2(_03236_),
    .A3(_03237_),
    .S0(net416),
    .S1(net414),
    .X(_03238_));
 sky130_fd_sc_hd__mux2i_4 _26497_ (.A0(_03233_),
    .A1(_03238_),
    .S(net413),
    .Y(_03239_));
 sky130_fd_sc_hd__mux4_2 _26498_ (.A0(\w[1][23] ),
    .A1(\w[5][23] ),
    .A2(\w[3][23] ),
    .A3(\w[7][23] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03240_));
 sky130_fd_sc_hd__mux4_2 _26499_ (.A0(\w[9][23] ),
    .A1(\w[13][23] ),
    .A2(\w[11][23] ),
    .A3(\w[15][23] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03241_));
 sky130_fd_sc_hd__mux4_2 _26500_ (.A0(\w[17][23] ),
    .A1(\w[21][23] ),
    .A2(\w[19][23] ),
    .A3(\w[23][23] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03242_));
 sky130_fd_sc_hd__mux4_2 _26501_ (.A0(\w[25][23] ),
    .A1(\w[29][23] ),
    .A2(\w[27][23] ),
    .A3(\w[31][23] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03243_));
 sky130_fd_sc_hd__mux4_2 _26502_ (.A0(_03240_),
    .A1(_03241_),
    .A2(_03242_),
    .A3(_03243_),
    .S0(\count2_2[3] ),
    .S1(net540),
    .X(_03244_));
 sky130_fd_sc_hd__mux4_2 _26503_ (.A0(\w[33][23] ),
    .A1(\w[37][23] ),
    .A2(\w[35][23] ),
    .A3(\w[39][23] ),
    .S0(net423),
    .S1(net428),
    .X(_03245_));
 sky130_fd_sc_hd__mux4_2 _26504_ (.A0(\w[41][23] ),
    .A1(\w[45][23] ),
    .A2(\w[43][23] ),
    .A3(\w[47][23] ),
    .S0(net423),
    .S1(net428),
    .X(_03246_));
 sky130_fd_sc_hd__mux4_2 _26505_ (.A0(\w[49][23] ),
    .A1(\w[53][23] ),
    .A2(\w[51][23] ),
    .A3(\w[55][23] ),
    .S0(net423),
    .S1(net428),
    .X(_03247_));
 sky130_fd_sc_hd__mux4_2 _26506_ (.A0(\w[57][23] ),
    .A1(\w[61][23] ),
    .A2(\w[59][23] ),
    .A3(\w[63][23] ),
    .S0(net423),
    .S1(net428),
    .X(_03248_));
 sky130_fd_sc_hd__mux4_2 _26507_ (.A0(_03245_),
    .A1(_03246_),
    .A2(_03247_),
    .A3(_03248_),
    .S0(net417),
    .S1(net414),
    .X(_03249_));
 sky130_fd_sc_hd__mux2i_4 _26508_ (.A0(_03244_),
    .A1(_03249_),
    .S(\count2_2[5] ),
    .Y(_03250_));
 sky130_fd_sc_hd__xnor2_1 _26509_ (.A(_03239_),
    .B(_03250_),
    .Y(_03251_));
 sky130_fd_sc_hd__xnor2_1 _26510_ (.A(_03086_),
    .B(_03251_),
    .Y(_11861_));
 sky130_fd_sc_hd__mux4_2 _26511_ (.A0(\w[0][22] ),
    .A1(\w[4][22] ),
    .A2(\w[2][22] ),
    .A3(\w[6][22] ),
    .S0(net500),
    .S1(net507),
    .X(_03252_));
 sky130_fd_sc_hd__mux4_2 _26512_ (.A0(\w[8][22] ),
    .A1(\w[12][22] ),
    .A2(\w[10][22] ),
    .A3(\w[14][22] ),
    .S0(net501),
    .S1(net507),
    .X(_03253_));
 sky130_fd_sc_hd__mux4_2 _26513_ (.A0(\w[16][22] ),
    .A1(\w[20][22] ),
    .A2(\w[18][22] ),
    .A3(\w[22][22] ),
    .S0(net501),
    .S1(net507),
    .X(_03254_));
 sky130_fd_sc_hd__mux4_2 _26514_ (.A0(\w[24][22] ),
    .A1(\w[28][22] ),
    .A2(\w[26][22] ),
    .A3(\w[30][22] ),
    .S0(net501),
    .S1(net507),
    .X(_03255_));
 sky130_fd_sc_hd__mux4_2 _26515_ (.A0(_03252_),
    .A1(_03253_),
    .A2(_03254_),
    .A3(_03255_),
    .S0(net497),
    .S1(net495),
    .X(_03256_));
 sky130_fd_sc_hd__mux4_2 _26516_ (.A0(\w[32][22] ),
    .A1(\w[36][22] ),
    .A2(\w[34][22] ),
    .A3(\w[38][22] ),
    .S0(net500),
    .S1(net507),
    .X(_03257_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_64 ();
 sky130_fd_sc_hd__mux4_2 _26518_ (.A0(\w[40][22] ),
    .A1(\w[44][22] ),
    .A2(\w[42][22] ),
    .A3(\w[46][22] ),
    .S0(net500),
    .S1(net507),
    .X(_03259_));
 sky130_fd_sc_hd__mux4_2 _26519_ (.A0(\w[48][22] ),
    .A1(\w[52][22] ),
    .A2(\w[50][22] ),
    .A3(\w[54][22] ),
    .S0(net500),
    .S1(net507),
    .X(_03260_));
 sky130_fd_sc_hd__mux4_2 _26520_ (.A0(\w[56][22] ),
    .A1(\w[60][22] ),
    .A2(\w[58][22] ),
    .A3(\w[62][22] ),
    .S0(net500),
    .S1(net507),
    .X(_03261_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_63 ();
 sky130_fd_sc_hd__mux4_2 _26522_ (.A0(_03257_),
    .A1(_03259_),
    .A2(_03260_),
    .A3(_03261_),
    .S0(net497),
    .S1(net495),
    .X(_03263_));
 sky130_fd_sc_hd__mux2i_4 _26523_ (.A0(_03256_),
    .A1(_03263_),
    .S(net492),
    .Y(_03264_));
 sky130_fd_sc_hd__mux4_2 _26524_ (.A0(\w[0][11] ),
    .A1(\w[4][11] ),
    .A2(\w[2][11] ),
    .A3(\w[6][11] ),
    .S0(net501),
    .S1(net507),
    .X(_03265_));
 sky130_fd_sc_hd__mux4_2 _26525_ (.A0(\w[8][11] ),
    .A1(\w[12][11] ),
    .A2(\w[10][11] ),
    .A3(\w[14][11] ),
    .S0(net498),
    .S1(net507),
    .X(_03266_));
 sky130_fd_sc_hd__mux4_2 _26526_ (.A0(\w[16][11] ),
    .A1(\w[20][11] ),
    .A2(\w[18][11] ),
    .A3(\w[22][11] ),
    .S0(net501),
    .S1(net507),
    .X(_03267_));
 sky130_fd_sc_hd__mux4_2 _26527_ (.A0(\w[24][11] ),
    .A1(\w[28][11] ),
    .A2(\w[26][11] ),
    .A3(\w[30][11] ),
    .S0(net501),
    .S1(net507),
    .X(_03268_));
 sky130_fd_sc_hd__mux4_2 _26528_ (.A0(_03265_),
    .A1(_03266_),
    .A2(_03267_),
    .A3(_03268_),
    .S0(net496),
    .S1(net494),
    .X(_03269_));
 sky130_fd_sc_hd__mux4_2 _26529_ (.A0(\w[32][11] ),
    .A1(\w[36][11] ),
    .A2(\w[34][11] ),
    .A3(\w[38][11] ),
    .S0(net504),
    .S1(net510),
    .X(_03270_));
 sky130_fd_sc_hd__mux4_2 _26530_ (.A0(\w[40][11] ),
    .A1(\w[44][11] ),
    .A2(\w[42][11] ),
    .A3(\w[46][11] ),
    .S0(net504),
    .S1(net510),
    .X(_03271_));
 sky130_fd_sc_hd__mux4_2 _26531_ (.A0(\w[48][11] ),
    .A1(\w[52][11] ),
    .A2(\w[50][11] ),
    .A3(\w[54][11] ),
    .S0(net504),
    .S1(net510),
    .X(_03272_));
 sky130_fd_sc_hd__mux4_2 _26532_ (.A0(\w[56][11] ),
    .A1(\w[60][11] ),
    .A2(\w[58][11] ),
    .A3(\w[62][11] ),
    .S0(net504),
    .S1(net510),
    .X(_03273_));
 sky130_fd_sc_hd__mux4_2 _26533_ (.A0(_03270_),
    .A1(_03271_),
    .A2(_03272_),
    .A3(_03273_),
    .S0(net497),
    .S1(net495),
    .X(_03274_));
 sky130_fd_sc_hd__mux2i_4 _26534_ (.A0(_03269_),
    .A1(_03274_),
    .S(net492),
    .Y(_03275_));
 sky130_fd_sc_hd__xnor2_1 _26535_ (.A(_03264_),
    .B(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__xnor2_2 _26536_ (.A(_02882_),
    .B(_03276_),
    .Y(_11860_));
 sky130_fd_sc_hd__mux4_2 _26537_ (.A0(\w[0][4] ),
    .A1(\w[4][4] ),
    .A2(\w[2][4] ),
    .A3(\w[6][4] ),
    .S0(net380),
    .S1(net388),
    .X(_03277_));
 sky130_fd_sc_hd__mux4_2 _26538_ (.A0(\w[8][4] ),
    .A1(\w[12][4] ),
    .A2(\w[10][4] ),
    .A3(\w[14][4] ),
    .S0(net380),
    .S1(net388),
    .X(_03278_));
 sky130_fd_sc_hd__mux4_2 _26539_ (.A0(\w[16][4] ),
    .A1(\w[20][4] ),
    .A2(\w[18][4] ),
    .A3(\w[22][4] ),
    .S0(net380),
    .S1(net388),
    .X(_03279_));
 sky130_fd_sc_hd__mux4_2 _26540_ (.A0(\w[24][4] ),
    .A1(\w[28][4] ),
    .A2(\w[26][4] ),
    .A3(\w[30][4] ),
    .S0(net380),
    .S1(net388),
    .X(_03280_));
 sky130_fd_sc_hd__mux4_2 _26541_ (.A0(_03277_),
    .A1(_03278_),
    .A2(_03279_),
    .A3(_03280_),
    .S0(net379),
    .S1(net376),
    .X(_03281_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_62 ();
 sky130_fd_sc_hd__mux4_2 _26543_ (.A0(\w[32][4] ),
    .A1(\w[36][4] ),
    .A2(\w[34][4] ),
    .A3(\w[38][4] ),
    .S0(net380),
    .S1(net388),
    .X(_03283_));
 sky130_fd_sc_hd__mux4_2 _26544_ (.A0(\w[40][4] ),
    .A1(\w[44][4] ),
    .A2(\w[42][4] ),
    .A3(\w[46][4] ),
    .S0(net380),
    .S1(net388),
    .X(_03284_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_61 ();
 sky130_fd_sc_hd__mux4_2 _26546_ (.A0(\w[48][4] ),
    .A1(\w[52][4] ),
    .A2(\w[50][4] ),
    .A3(\w[54][4] ),
    .S0(net380),
    .S1(net388),
    .X(_03286_));
 sky130_fd_sc_hd__mux4_2 _26547_ (.A0(\w[56][4] ),
    .A1(\w[60][4] ),
    .A2(\w[58][4] ),
    .A3(\w[62][4] ),
    .S0(net380),
    .S1(net388),
    .X(_03287_));
 sky130_fd_sc_hd__mux4_2 _26548_ (.A0(_03283_),
    .A1(_03284_),
    .A2(_03286_),
    .A3(_03287_),
    .S0(net379),
    .S1(net376),
    .X(_03288_));
 sky130_fd_sc_hd__mux2i_4 _26549_ (.A0(_03281_),
    .A1(_03288_),
    .S(net373),
    .Y(_11859_));
 sky130_fd_sc_hd__mux4_2 _26550_ (.A0(\w[1][4] ),
    .A1(\w[5][4] ),
    .A2(\w[3][4] ),
    .A3(\w[7][4] ),
    .S0(net460),
    .S1(net470),
    .X(_03289_));
 sky130_fd_sc_hd__mux4_2 _26551_ (.A0(\w[9][4] ),
    .A1(\w[13][4] ),
    .A2(\w[11][4] ),
    .A3(\w[15][4] ),
    .S0(net460),
    .S1(net470),
    .X(_03290_));
 sky130_fd_sc_hd__mux4_2 _26552_ (.A0(\w[17][4] ),
    .A1(\w[21][4] ),
    .A2(\w[19][4] ),
    .A3(\w[23][4] ),
    .S0(net460),
    .S1(net470),
    .X(_03291_));
 sky130_fd_sc_hd__mux4_2 _26553_ (.A0(\w[25][4] ),
    .A1(\w[29][4] ),
    .A2(\w[27][4] ),
    .A3(\w[31][4] ),
    .S0(net460),
    .S1(net470),
    .X(_03292_));
 sky130_fd_sc_hd__mux4_2 _26554_ (.A0(_03289_),
    .A1(_03290_),
    .A2(_03291_),
    .A3(_03292_),
    .S0(net456),
    .S1(net454),
    .X(_03293_));
 sky130_fd_sc_hd__mux4_2 _26555_ (.A0(\w[33][4] ),
    .A1(\w[37][4] ),
    .A2(\w[35][4] ),
    .A3(\w[39][4] ),
    .S0(net460),
    .S1(net468),
    .X(_03294_));
 sky130_fd_sc_hd__mux4_2 _26556_ (.A0(\w[41][4] ),
    .A1(\w[45][4] ),
    .A2(\w[43][4] ),
    .A3(\w[47][4] ),
    .S0(net460),
    .S1(net468),
    .X(_03295_));
 sky130_fd_sc_hd__mux4_2 _26557_ (.A0(\w[49][4] ),
    .A1(\w[53][4] ),
    .A2(\w[51][4] ),
    .A3(\w[55][4] ),
    .S0(net460),
    .S1(net468),
    .X(_03296_));
 sky130_fd_sc_hd__mux4_2 _26558_ (.A0(\w[57][4] ),
    .A1(\w[61][4] ),
    .A2(\w[59][4] ),
    .A3(\w[63][4] ),
    .S0(net460),
    .S1(net469),
    .X(_03297_));
 sky130_fd_sc_hd__mux4_2 _26559_ (.A0(_03294_),
    .A1(_03295_),
    .A2(_03296_),
    .A3(_03297_),
    .S0(net456),
    .S1(net454),
    .X(_03298_));
 sky130_fd_sc_hd__mux2i_2 _26560_ (.A0(_03293_),
    .A1(_03298_),
    .S(net453),
    .Y(_11864_));
 sky130_fd_sc_hd__mux4_2 _26561_ (.A0(\w[1][15] ),
    .A1(\w[5][15] ),
    .A2(\w[3][15] ),
    .A3(\w[7][15] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03299_));
 sky130_fd_sc_hd__mux4_2 _26562_ (.A0(\w[9][15] ),
    .A1(\w[13][15] ),
    .A2(\w[11][15] ),
    .A3(\w[15][15] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03300_));
 sky130_fd_sc_hd__mux4_2 _26563_ (.A0(\w[17][15] ),
    .A1(\w[21][15] ),
    .A2(\w[19][15] ),
    .A3(\w[23][15] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03301_));
 sky130_fd_sc_hd__mux4_2 _26564_ (.A0(\w[25][15] ),
    .A1(\w[29][15] ),
    .A2(\w[27][15] ),
    .A3(\w[31][15] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03302_));
 sky130_fd_sc_hd__mux4_2 _26565_ (.A0(_03299_),
    .A1(_03300_),
    .A2(_03301_),
    .A3(_03302_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[4] ),
    .X(_03303_));
 sky130_fd_sc_hd__mux4_2 _26566_ (.A0(\w[33][15] ),
    .A1(\w[37][15] ),
    .A2(\w[35][15] ),
    .A3(\w[39][15] ),
    .S0(net425),
    .S1(net430),
    .X(_03304_));
 sky130_fd_sc_hd__mux4_2 _26567_ (.A0(\w[41][15] ),
    .A1(\w[45][15] ),
    .A2(\w[43][15] ),
    .A3(\w[47][15] ),
    .S0(net425),
    .S1(net430),
    .X(_03305_));
 sky130_fd_sc_hd__mux4_2 _26568_ (.A0(\w[49][15] ),
    .A1(\w[53][15] ),
    .A2(\w[51][15] ),
    .A3(\w[55][15] ),
    .S0(net425),
    .S1(net430),
    .X(_03306_));
 sky130_fd_sc_hd__mux4_2 _26569_ (.A0(\w[57][15] ),
    .A1(\w[61][15] ),
    .A2(\w[59][15] ),
    .A3(\w[63][15] ),
    .S0(net425),
    .S1(net430),
    .X(_03307_));
 sky130_fd_sc_hd__mux4_2 _26570_ (.A0(_03304_),
    .A1(_03305_),
    .A2(_03306_),
    .A3(_03307_),
    .S0(net418),
    .S1(\count2_2[4] ),
    .X(_03308_));
 sky130_fd_sc_hd__mux2i_4 _26571_ (.A0(_03303_),
    .A1(_03308_),
    .S(\count2_2[5] ),
    .Y(_03309_));
 sky130_fd_sc_hd__mux4_2 _26572_ (.A0(\w[1][24] ),
    .A1(\w[5][24] ),
    .A2(\w[3][24] ),
    .A3(\w[7][24] ),
    .S0(net422),
    .S1(net429),
    .X(_03310_));
 sky130_fd_sc_hd__mux4_2 _26573_ (.A0(\w[9][24] ),
    .A1(\w[13][24] ),
    .A2(\w[11][24] ),
    .A3(\w[15][24] ),
    .S0(net422),
    .S1(net429),
    .X(_03311_));
 sky130_fd_sc_hd__mux4_2 _26574_ (.A0(\w[17][24] ),
    .A1(\w[21][24] ),
    .A2(\w[19][24] ),
    .A3(\w[23][24] ),
    .S0(net422),
    .S1(net429),
    .X(_03312_));
 sky130_fd_sc_hd__mux4_2 _26575_ (.A0(\w[25][24] ),
    .A1(\w[29][24] ),
    .A2(\w[27][24] ),
    .A3(\w[31][24] ),
    .S0(net422),
    .S1(net429),
    .X(_03313_));
 sky130_fd_sc_hd__mux4_2 _26576_ (.A0(_03310_),
    .A1(_03311_),
    .A2(_03312_),
    .A3(_03313_),
    .S0(net416),
    .S1(net414),
    .X(_03314_));
 sky130_fd_sc_hd__mux4_2 _26577_ (.A0(\w[33][24] ),
    .A1(\w[37][24] ),
    .A2(\w[35][24] ),
    .A3(\w[39][24] ),
    .S0(net423),
    .S1(net428),
    .X(_03315_));
 sky130_fd_sc_hd__mux4_2 _26578_ (.A0(\w[41][24] ),
    .A1(\w[45][24] ),
    .A2(\w[43][24] ),
    .A3(\w[47][24] ),
    .S0(net421),
    .S1(net428),
    .X(_03316_));
 sky130_fd_sc_hd__mux4_2 _26579_ (.A0(\w[49][24] ),
    .A1(\w[53][24] ),
    .A2(\w[51][24] ),
    .A3(\w[55][24] ),
    .S0(net423),
    .S1(net428),
    .X(_03317_));
 sky130_fd_sc_hd__mux4_2 _26580_ (.A0(\w[57][24] ),
    .A1(\w[61][24] ),
    .A2(\w[59][24] ),
    .A3(\w[63][24] ),
    .S0(net421),
    .S1(net428),
    .X(_03318_));
 sky130_fd_sc_hd__mux4_2 _26581_ (.A0(_03315_),
    .A1(_03316_),
    .A2(_03317_),
    .A3(_03318_),
    .S0(net417),
    .S1(net414),
    .X(_03319_));
 sky130_fd_sc_hd__mux2i_4 _26582_ (.A0(_03314_),
    .A1(_03319_),
    .S(net539),
    .Y(_03320_));
 sky130_fd_sc_hd__xnor2_1 _26583_ (.A(_03309_),
    .B(_03320_),
    .Y(_03321_));
 sky130_fd_sc_hd__xnor2_1 _26584_ (.A(_03168_),
    .B(_03321_),
    .Y(_11869_));
 sky130_fd_sc_hd__mux4_2 _26585_ (.A0(\w[0][23] ),
    .A1(\w[4][23] ),
    .A2(\w[2][23] ),
    .A3(\w[6][23] ),
    .S0(net498),
    .S1(net511),
    .X(_03322_));
 sky130_fd_sc_hd__mux4_2 _26586_ (.A0(\w[8][23] ),
    .A1(\w[12][23] ),
    .A2(\w[10][23] ),
    .A3(\w[14][23] ),
    .S0(net498),
    .S1(net511),
    .X(_03323_));
 sky130_fd_sc_hd__mux4_2 _26587_ (.A0(\w[16][23] ),
    .A1(\w[20][23] ),
    .A2(\w[18][23] ),
    .A3(\w[22][23] ),
    .S0(net498),
    .S1(net511),
    .X(_03324_));
 sky130_fd_sc_hd__mux4_2 _26588_ (.A0(\w[24][23] ),
    .A1(\w[28][23] ),
    .A2(\w[26][23] ),
    .A3(\w[30][23] ),
    .S0(net498),
    .S1(net511),
    .X(_03325_));
 sky130_fd_sc_hd__mux4_2 _26589_ (.A0(_03322_),
    .A1(_03323_),
    .A2(_03324_),
    .A3(_03325_),
    .S0(net496),
    .S1(net494),
    .X(_03326_));
 sky130_fd_sc_hd__mux4_2 _26590_ (.A0(\w[32][23] ),
    .A1(\w[36][23] ),
    .A2(\w[34][23] ),
    .A3(\w[38][23] ),
    .S0(net503),
    .S1(net509),
    .X(_03327_));
 sky130_fd_sc_hd__mux4_2 _26591_ (.A0(\w[40][23] ),
    .A1(\w[44][23] ),
    .A2(\w[42][23] ),
    .A3(\w[46][23] ),
    .S0(net503),
    .S1(net509),
    .X(_03328_));
 sky130_fd_sc_hd__mux4_2 _26592_ (.A0(\w[48][23] ),
    .A1(\w[52][23] ),
    .A2(\w[50][23] ),
    .A3(\w[54][23] ),
    .S0(net503),
    .S1(net509),
    .X(_03329_));
 sky130_fd_sc_hd__mux4_2 _26593_ (.A0(\w[56][23] ),
    .A1(\w[60][23] ),
    .A2(\w[58][23] ),
    .A3(\w[62][23] ),
    .S0(net503),
    .S1(net509),
    .X(_03330_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_60 ();
 sky130_fd_sc_hd__mux4_2 _26595_ (.A0(_03327_),
    .A1(_03328_),
    .A2(_03329_),
    .A3(_03330_),
    .S0(\count15_2[3] ),
    .S1(net494),
    .X(_03332_));
 sky130_fd_sc_hd__mux2i_4 _26596_ (.A0(_03326_),
    .A1(_03332_),
    .S(net493),
    .Y(_03333_));
 sky130_fd_sc_hd__mux4_2 _26597_ (.A0(\w[0][12] ),
    .A1(\w[4][12] ),
    .A2(\w[2][12] ),
    .A3(\w[6][12] ),
    .S0(net498),
    .S1(net511),
    .X(_03334_));
 sky130_fd_sc_hd__mux4_2 _26598_ (.A0(\w[8][12] ),
    .A1(\w[12][12] ),
    .A2(\w[10][12] ),
    .A3(\w[14][12] ),
    .S0(net498),
    .S1(net511),
    .X(_03335_));
 sky130_fd_sc_hd__mux4_2 _26599_ (.A0(\w[16][12] ),
    .A1(\w[20][12] ),
    .A2(\w[18][12] ),
    .A3(\w[22][12] ),
    .S0(net498),
    .S1(net511),
    .X(_03336_));
 sky130_fd_sc_hd__mux4_2 _26600_ (.A0(\w[24][12] ),
    .A1(\w[28][12] ),
    .A2(\w[26][12] ),
    .A3(\w[30][12] ),
    .S0(net498),
    .S1(net511),
    .X(_03337_));
 sky130_fd_sc_hd__mux4_2 _26601_ (.A0(_03334_),
    .A1(_03335_),
    .A2(_03336_),
    .A3(_03337_),
    .S0(net496),
    .S1(net547),
    .X(_03338_));
 sky130_fd_sc_hd__mux4_2 _26602_ (.A0(\w[32][12] ),
    .A1(\w[36][12] ),
    .A2(\w[34][12] ),
    .A3(\w[38][12] ),
    .S0(net505),
    .S1(net511),
    .X(_03339_));
 sky130_fd_sc_hd__mux4_2 _26603_ (.A0(\w[40][12] ),
    .A1(\w[44][12] ),
    .A2(\w[42][12] ),
    .A3(\w[46][12] ),
    .S0(net505),
    .S1(net511),
    .X(_03340_));
 sky130_fd_sc_hd__mux4_2 _26604_ (.A0(\w[48][12] ),
    .A1(\w[52][12] ),
    .A2(\w[50][12] ),
    .A3(\w[54][12] ),
    .S0(net505),
    .S1(net511),
    .X(_03341_));
 sky130_fd_sc_hd__mux4_2 _26605_ (.A0(\w[56][12] ),
    .A1(\w[60][12] ),
    .A2(\w[58][12] ),
    .A3(\w[62][12] ),
    .S0(net505),
    .S1(net511),
    .X(_03342_));
 sky130_fd_sc_hd__mux4_2 _26606_ (.A0(_03339_),
    .A1(_03340_),
    .A2(_03341_),
    .A3(_03342_),
    .S0(\count15_2[3] ),
    .S1(net494),
    .X(_03343_));
 sky130_fd_sc_hd__mux2i_4 _26607_ (.A0(_03338_),
    .A1(_03343_),
    .S(net493),
    .Y(_03344_));
 sky130_fd_sc_hd__xnor2_1 _26608_ (.A(_03333_),
    .B(_03344_),
    .Y(_03345_));
 sky130_fd_sc_hd__xnor2_1 _26609_ (.A(_02994_),
    .B(_03345_),
    .Y(_11868_));
 sky130_fd_sc_hd__mux4_2 _26610_ (.A0(\w[0][5] ),
    .A1(\w[4][5] ),
    .A2(\w[2][5] ),
    .A3(\w[6][5] ),
    .S0(net380),
    .S1(net388),
    .X(_03346_));
 sky130_fd_sc_hd__mux4_2 _26611_ (.A0(\w[8][5] ),
    .A1(\w[12][5] ),
    .A2(\w[10][5] ),
    .A3(\w[14][5] ),
    .S0(net380),
    .S1(net388),
    .X(_03347_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_59 ();
 sky130_fd_sc_hd__mux4_2 _26613_ (.A0(\w[16][5] ),
    .A1(\w[20][5] ),
    .A2(\w[18][5] ),
    .A3(\w[22][5] ),
    .S0(net380),
    .S1(net388),
    .X(_03349_));
 sky130_fd_sc_hd__mux4_2 _26614_ (.A0(\w[24][5] ),
    .A1(\w[28][5] ),
    .A2(\w[26][5] ),
    .A3(\w[30][5] ),
    .S0(net380),
    .S1(net388),
    .X(_03350_));
 sky130_fd_sc_hd__mux4_2 _26615_ (.A0(_03346_),
    .A1(_03347_),
    .A2(_03349_),
    .A3(_03350_),
    .S0(\count7_2[3] ),
    .S1(net376),
    .X(_03351_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_58 ();
 sky130_fd_sc_hd__mux4_2 _26617_ (.A0(\w[32][5] ),
    .A1(\w[36][5] ),
    .A2(\w[34][5] ),
    .A3(\w[38][5] ),
    .S0(net380),
    .S1(net388),
    .X(_03353_));
 sky130_fd_sc_hd__mux4_2 _26618_ (.A0(\w[40][5] ),
    .A1(\w[44][5] ),
    .A2(\w[42][5] ),
    .A3(\w[46][5] ),
    .S0(net380),
    .S1(net388),
    .X(_03354_));
 sky130_fd_sc_hd__mux4_2 _26619_ (.A0(\w[48][5] ),
    .A1(\w[52][5] ),
    .A2(\w[50][5] ),
    .A3(\w[54][5] ),
    .S0(net380),
    .S1(net388),
    .X(_03355_));
 sky130_fd_sc_hd__mux4_2 _26620_ (.A0(\w[56][5] ),
    .A1(\w[60][5] ),
    .A2(\w[58][5] ),
    .A3(\w[62][5] ),
    .S0(net387),
    .S1(net388),
    .X(_03356_));
 sky130_fd_sc_hd__mux4_2 _26621_ (.A0(_03353_),
    .A1(_03354_),
    .A2(_03355_),
    .A3(_03356_),
    .S0(net379),
    .S1(net376),
    .X(_03357_));
 sky130_fd_sc_hd__mux2i_4 _26622_ (.A0(_03351_),
    .A1(_03357_),
    .S(net373),
    .Y(_11867_));
 sky130_fd_sc_hd__mux4_2 _26623_ (.A0(\w[1][5] ),
    .A1(\w[5][5] ),
    .A2(\w[3][5] ),
    .A3(\w[7][5] ),
    .S0(net459),
    .S1(net544),
    .X(_03358_));
 sky130_fd_sc_hd__mux4_2 _26624_ (.A0(\w[9][5] ),
    .A1(\w[13][5] ),
    .A2(\w[11][5] ),
    .A3(\w[15][5] ),
    .S0(net459),
    .S1(net544),
    .X(_03359_));
 sky130_fd_sc_hd__mux4_2 _26625_ (.A0(\w[17][5] ),
    .A1(\w[21][5] ),
    .A2(\w[19][5] ),
    .A3(\w[23][5] ),
    .S0(net459),
    .S1(net544),
    .X(_03360_));
 sky130_fd_sc_hd__mux4_2 _26626_ (.A0(\w[25][5] ),
    .A1(\w[29][5] ),
    .A2(\w[27][5] ),
    .A3(\w[31][5] ),
    .S0(net461),
    .S1(net544),
    .X(_03361_));
 sky130_fd_sc_hd__mux4_2 _26627_ (.A0(_03358_),
    .A1(_03359_),
    .A2(_03360_),
    .A3(_03361_),
    .S0(net456),
    .S1(net454),
    .X(_03362_));
 sky130_fd_sc_hd__mux4_2 _26628_ (.A0(\w[33][5] ),
    .A1(\w[37][5] ),
    .A2(\w[35][5] ),
    .A3(\w[39][5] ),
    .S0(net461),
    .S1(net544),
    .X(_03363_));
 sky130_fd_sc_hd__mux4_2 _26629_ (.A0(\w[41][5] ),
    .A1(\w[45][5] ),
    .A2(\w[43][5] ),
    .A3(\w[47][5] ),
    .S0(net461),
    .S1(net544),
    .X(_03364_));
 sky130_fd_sc_hd__mux4_2 _26630_ (.A0(\w[49][5] ),
    .A1(\w[53][5] ),
    .A2(\w[51][5] ),
    .A3(\w[55][5] ),
    .S0(net461),
    .S1(net544),
    .X(_03365_));
 sky130_fd_sc_hd__mux4_2 _26631_ (.A0(\w[57][5] ),
    .A1(\w[61][5] ),
    .A2(\w[59][5] ),
    .A3(\w[63][5] ),
    .S0(net461),
    .S1(net544),
    .X(_03366_));
 sky130_fd_sc_hd__mux4_2 _26632_ (.A0(_03363_),
    .A1(_03364_),
    .A2(_03365_),
    .A3(_03366_),
    .S0(net456),
    .S1(net543),
    .X(_03367_));
 sky130_fd_sc_hd__mux2i_4 _26633_ (.A0(_03362_),
    .A1(_03367_),
    .S(net453),
    .Y(_11872_));
 sky130_fd_sc_hd__mux4_2 _26634_ (.A0(\w[1][16] ),
    .A1(\w[5][16] ),
    .A2(\w[3][16] ),
    .A3(\w[7][16] ),
    .S0(net423),
    .S1(net427),
    .X(_03368_));
 sky130_fd_sc_hd__mux4_2 _26635_ (.A0(\w[9][16] ),
    .A1(\w[13][16] ),
    .A2(\w[11][16] ),
    .A3(\w[15][16] ),
    .S0(net423),
    .S1(net427),
    .X(_03369_));
 sky130_fd_sc_hd__mux4_2 _26636_ (.A0(\w[17][16] ),
    .A1(\w[21][16] ),
    .A2(\w[19][16] ),
    .A3(\w[23][16] ),
    .S0(net423),
    .S1(net427),
    .X(_03370_));
 sky130_fd_sc_hd__mux4_2 _26637_ (.A0(\w[25][16] ),
    .A1(\w[29][16] ),
    .A2(\w[27][16] ),
    .A3(\w[31][16] ),
    .S0(net423),
    .S1(net427),
    .X(_03371_));
 sky130_fd_sc_hd__mux4_2 _26638_ (.A0(_03368_),
    .A1(_03369_),
    .A2(_03370_),
    .A3(_03371_),
    .S0(net416),
    .S1(net414),
    .X(_03372_));
 sky130_fd_sc_hd__mux4_2 _26639_ (.A0(\w[33][16] ),
    .A1(\w[37][16] ),
    .A2(\w[35][16] ),
    .A3(\w[39][16] ),
    .S0(net421),
    .S1(net428),
    .X(_03373_));
 sky130_fd_sc_hd__mux4_2 _26640_ (.A0(\w[41][16] ),
    .A1(\w[45][16] ),
    .A2(\w[43][16] ),
    .A3(\w[47][16] ),
    .S0(net419),
    .S1(net426),
    .X(_03374_));
 sky130_fd_sc_hd__mux4_2 _26641_ (.A0(\w[49][16] ),
    .A1(\w[53][16] ),
    .A2(\w[51][16] ),
    .A3(\w[55][16] ),
    .S0(net421),
    .S1(net428),
    .X(_03375_));
 sky130_fd_sc_hd__mux4_2 _26642_ (.A0(\w[57][16] ),
    .A1(\w[61][16] ),
    .A2(\w[59][16] ),
    .A3(\w[63][16] ),
    .S0(net421),
    .S1(net428),
    .X(_03376_));
 sky130_fd_sc_hd__mux4_2 _26643_ (.A0(_03373_),
    .A1(_03374_),
    .A2(_03375_),
    .A3(_03376_),
    .S0(net417),
    .S1(net414),
    .X(_03377_));
 sky130_fd_sc_hd__mux2i_4 _26644_ (.A0(_03372_),
    .A1(_03377_),
    .S(net539),
    .Y(_03378_));
 sky130_fd_sc_hd__mux4_2 _26645_ (.A0(\w[1][25] ),
    .A1(\w[5][25] ),
    .A2(\w[3][25] ),
    .A3(\w[7][25] ),
    .S0(net420),
    .S1(net427),
    .X(_03379_));
 sky130_fd_sc_hd__mux4_2 _26646_ (.A0(\w[9][25] ),
    .A1(\w[13][25] ),
    .A2(\w[11][25] ),
    .A3(\w[15][25] ),
    .S0(net420),
    .S1(net427),
    .X(_03380_));
 sky130_fd_sc_hd__mux4_2 _26647_ (.A0(\w[17][25] ),
    .A1(\w[21][25] ),
    .A2(\w[19][25] ),
    .A3(\w[23][25] ),
    .S0(net420),
    .S1(net427),
    .X(_03381_));
 sky130_fd_sc_hd__mux4_2 _26648_ (.A0(\w[25][25] ),
    .A1(\w[29][25] ),
    .A2(\w[27][25] ),
    .A3(\w[31][25] ),
    .S0(net420),
    .S1(net427),
    .X(_03382_));
 sky130_fd_sc_hd__mux4_2 _26649_ (.A0(_03379_),
    .A1(_03380_),
    .A2(_03381_),
    .A3(_03382_),
    .S0(net416),
    .S1(net415),
    .X(_03383_));
 sky130_fd_sc_hd__mux4_2 _26650_ (.A0(\w[33][25] ),
    .A1(\w[37][25] ),
    .A2(\w[35][25] ),
    .A3(\w[39][25] ),
    .S0(net420),
    .S1(net427),
    .X(_03384_));
 sky130_fd_sc_hd__mux4_2 _26651_ (.A0(\w[41][25] ),
    .A1(\w[45][25] ),
    .A2(\w[43][25] ),
    .A3(\w[47][25] ),
    .S0(net420),
    .S1(net427),
    .X(_03385_));
 sky130_fd_sc_hd__mux4_2 _26652_ (.A0(\w[49][25] ),
    .A1(\w[53][25] ),
    .A2(\w[51][25] ),
    .A3(\w[55][25] ),
    .S0(net420),
    .S1(net427),
    .X(_03386_));
 sky130_fd_sc_hd__mux4_2 _26653_ (.A0(\w[57][25] ),
    .A1(\w[61][25] ),
    .A2(\w[59][25] ),
    .A3(\w[63][25] ),
    .S0(net420),
    .S1(net427),
    .X(_03387_));
 sky130_fd_sc_hd__mux4_2 _26654_ (.A0(_03384_),
    .A1(_03385_),
    .A2(_03386_),
    .A3(_03387_),
    .S0(net417),
    .S1(net415),
    .X(_03388_));
 sky130_fd_sc_hd__mux2i_4 _26655_ (.A0(_03383_),
    .A1(_03388_),
    .S(net413),
    .Y(_03389_));
 sky130_fd_sc_hd__xnor2_1 _26656_ (.A(_03378_),
    .B(_03389_),
    .Y(_03390_));
 sky130_fd_sc_hd__xnor2_1 _26657_ (.A(_03250_),
    .B(_03390_),
    .Y(_11877_));
 sky130_fd_sc_hd__mux4_2 _26658_ (.A0(\w[0][13] ),
    .A1(\w[4][13] ),
    .A2(\w[2][13] ),
    .A3(\w[6][13] ),
    .S0(net503),
    .S1(net509),
    .X(_03391_));
 sky130_fd_sc_hd__mux4_2 _26659_ (.A0(\w[8][13] ),
    .A1(\w[12][13] ),
    .A2(\w[10][13] ),
    .A3(\w[14][13] ),
    .S0(net503),
    .S1(net509),
    .X(_03392_));
 sky130_fd_sc_hd__mux4_2 _26660_ (.A0(\w[16][13] ),
    .A1(\w[20][13] ),
    .A2(\w[18][13] ),
    .A3(\w[22][13] ),
    .S0(net503),
    .S1(net509),
    .X(_03393_));
 sky130_fd_sc_hd__mux4_2 _26661_ (.A0(\w[24][13] ),
    .A1(\w[28][13] ),
    .A2(\w[26][13] ),
    .A3(\w[30][13] ),
    .S0(net503),
    .S1(net509),
    .X(_03394_));
 sky130_fd_sc_hd__mux4_2 _26662_ (.A0(_03391_),
    .A1(_03392_),
    .A2(_03393_),
    .A3(_03394_),
    .S0(net496),
    .S1(net494),
    .X(_03395_));
 sky130_fd_sc_hd__mux4_2 _26663_ (.A0(\w[32][13] ),
    .A1(\w[36][13] ),
    .A2(\w[34][13] ),
    .A3(\w[38][13] ),
    .S0(net504),
    .S1(net510),
    .X(_03396_));
 sky130_fd_sc_hd__mux4_2 _26664_ (.A0(\w[40][13] ),
    .A1(\w[44][13] ),
    .A2(\w[42][13] ),
    .A3(\w[46][13] ),
    .S0(net504),
    .S1(net510),
    .X(_03397_));
 sky130_fd_sc_hd__mux4_2 _26665_ (.A0(\w[48][13] ),
    .A1(\w[52][13] ),
    .A2(\w[50][13] ),
    .A3(\w[54][13] ),
    .S0(net505),
    .S1(net511),
    .X(_03398_));
 sky130_fd_sc_hd__mux4_2 _26666_ (.A0(\w[56][13] ),
    .A1(\w[60][13] ),
    .A2(\w[58][13] ),
    .A3(\w[62][13] ),
    .S0(net505),
    .S1(net511),
    .X(_03399_));
 sky130_fd_sc_hd__mux4_2 _26667_ (.A0(_03396_),
    .A1(_03397_),
    .A2(_03398_),
    .A3(_03399_),
    .S0(net497),
    .S1(\count15_2[4] ),
    .X(_03400_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_57 ();
 sky130_fd_sc_hd__mux2i_4 _26669_ (.A0(_03395_),
    .A1(_03400_),
    .S(net493),
    .Y(_03402_));
 sky130_fd_sc_hd__mux4_2 _26670_ (.A0(\w[0][24] ),
    .A1(\w[4][24] ),
    .A2(\w[2][24] ),
    .A3(\w[6][24] ),
    .S0(net500),
    .S1(net507),
    .X(_03403_));
 sky130_fd_sc_hd__mux4_2 _26671_ (.A0(\w[8][24] ),
    .A1(\w[12][24] ),
    .A2(\w[10][24] ),
    .A3(\w[14][24] ),
    .S0(net500),
    .S1(net507),
    .X(_03404_));
 sky130_fd_sc_hd__mux4_2 _26672_ (.A0(\w[16][24] ),
    .A1(\w[20][24] ),
    .A2(\w[18][24] ),
    .A3(\w[22][24] ),
    .S0(net500),
    .S1(net507),
    .X(_03405_));
 sky130_fd_sc_hd__mux4_2 _26673_ (.A0(\w[24][24] ),
    .A1(\w[28][24] ),
    .A2(\w[26][24] ),
    .A3(\w[30][24] ),
    .S0(net500),
    .S1(net507),
    .X(_03406_));
 sky130_fd_sc_hd__mux4_2 _26674_ (.A0(_03403_),
    .A1(_03404_),
    .A2(_03405_),
    .A3(_03406_),
    .S0(net497),
    .S1(net495),
    .X(_03407_));
 sky130_fd_sc_hd__mux4_2 _26675_ (.A0(\w[32][24] ),
    .A1(\w[36][24] ),
    .A2(\w[34][24] ),
    .A3(\w[38][24] ),
    .S0(net501),
    .S1(net507),
    .X(_03408_));
 sky130_fd_sc_hd__mux4_2 _26676_ (.A0(\w[40][24] ),
    .A1(\w[44][24] ),
    .A2(\w[42][24] ),
    .A3(\w[46][24] ),
    .S0(net500),
    .S1(net507),
    .X(_03409_));
 sky130_fd_sc_hd__mux4_2 _26677_ (.A0(\w[48][24] ),
    .A1(\w[52][24] ),
    .A2(\w[50][24] ),
    .A3(\w[54][24] ),
    .S0(net501),
    .S1(net507),
    .X(_03410_));
 sky130_fd_sc_hd__mux4_2 _26678_ (.A0(\w[56][24] ),
    .A1(\w[60][24] ),
    .A2(\w[58][24] ),
    .A3(\w[62][24] ),
    .S0(net501),
    .S1(net507),
    .X(_03411_));
 sky130_fd_sc_hd__mux4_2 _26679_ (.A0(_03408_),
    .A1(_03409_),
    .A2(_03410_),
    .A3(_03411_),
    .S0(net497),
    .S1(net495),
    .X(_03412_));
 sky130_fd_sc_hd__mux2i_4 _26680_ (.A0(_03407_),
    .A1(_03412_),
    .S(net492),
    .Y(_03413_));
 sky130_fd_sc_hd__xnor2_1 _26681_ (.A(_03402_),
    .B(_03413_),
    .Y(_03414_));
 sky130_fd_sc_hd__xnor2_1 _26682_ (.A(_03120_),
    .B(_03414_),
    .Y(_11876_));
 sky130_fd_sc_hd__mux4_2 _26683_ (.A0(\w[0][6] ),
    .A1(\w[4][6] ),
    .A2(\w[2][6] ),
    .A3(\w[6][6] ),
    .S0(net387),
    .S1(net388),
    .X(_03415_));
 sky130_fd_sc_hd__mux4_2 _26684_ (.A0(\w[8][6] ),
    .A1(\w[12][6] ),
    .A2(\w[10][6] ),
    .A3(\w[14][6] ),
    .S0(net387),
    .S1(net388),
    .X(_03416_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_56 ();
 sky130_fd_sc_hd__mux4_2 _26686_ (.A0(\w[16][6] ),
    .A1(\w[20][6] ),
    .A2(\w[18][6] ),
    .A3(\w[22][6] ),
    .S0(net387),
    .S1(net388),
    .X(_03418_));
 sky130_fd_sc_hd__mux4_2 _26687_ (.A0(\w[24][6] ),
    .A1(\w[28][6] ),
    .A2(\w[26][6] ),
    .A3(\w[30][6] ),
    .S0(net387),
    .S1(net388),
    .X(_03419_));
 sky130_fd_sc_hd__mux4_2 _26688_ (.A0(_03415_),
    .A1(_03416_),
    .A2(_03418_),
    .A3(_03419_),
    .S0(\count7_2[3] ),
    .S1(net376),
    .X(_03420_));
 sky130_fd_sc_hd__mux4_2 _26689_ (.A0(\w[32][6] ),
    .A1(\w[36][6] ),
    .A2(\w[34][6] ),
    .A3(\w[38][6] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_03421_));
 sky130_fd_sc_hd__mux4_2 _26690_ (.A0(\w[40][6] ),
    .A1(\w[44][6] ),
    .A2(\w[42][6] ),
    .A3(\w[46][6] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_03422_));
 sky130_fd_sc_hd__mux4_2 _26691_ (.A0(\w[48][6] ),
    .A1(\w[52][6] ),
    .A2(\w[50][6] ),
    .A3(\w[54][6] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_03423_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_55 ();
 sky130_fd_sc_hd__mux4_2 _26693_ (.A0(\w[56][6] ),
    .A1(\w[60][6] ),
    .A2(\w[58][6] ),
    .A3(\w[62][6] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_03425_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_54 ();
 sky130_fd_sc_hd__mux4_2 _26695_ (.A0(_03421_),
    .A1(_03422_),
    .A2(_03423_),
    .A3(_03425_),
    .S0(net379),
    .S1(net376),
    .X(_03427_));
 sky130_fd_sc_hd__mux2i_4 _26696_ (.A0(_03420_),
    .A1(_03427_),
    .S(net374),
    .Y(_11875_));
 sky130_fd_sc_hd__mux4_2 _26697_ (.A0(\w[1][6] ),
    .A1(\w[5][6] ),
    .A2(\w[3][6] ),
    .A3(\w[7][6] ),
    .S0(net464),
    .S1(net468),
    .X(_03428_));
 sky130_fd_sc_hd__mux4_2 _26698_ (.A0(\w[9][6] ),
    .A1(\w[13][6] ),
    .A2(\w[11][6] ),
    .A3(\w[15][6] ),
    .S0(net464),
    .S1(net468),
    .X(_03429_));
 sky130_fd_sc_hd__mux4_2 _26699_ (.A0(\w[17][6] ),
    .A1(\w[21][6] ),
    .A2(\w[19][6] ),
    .A3(\w[23][6] ),
    .S0(net464),
    .S1(net468),
    .X(_03430_));
 sky130_fd_sc_hd__mux4_2 _26700_ (.A0(\w[25][6] ),
    .A1(\w[29][6] ),
    .A2(\w[27][6] ),
    .A3(\w[31][6] ),
    .S0(net464),
    .S1(net468),
    .X(_03431_));
 sky130_fd_sc_hd__mux4_2 _26701_ (.A0(_03428_),
    .A1(_03429_),
    .A2(_03430_),
    .A3(_03431_),
    .S0(\count16_2[3] ),
    .S1(net454),
    .X(_03432_));
 sky130_fd_sc_hd__mux4_2 _26702_ (.A0(\w[33][6] ),
    .A1(\w[37][6] ),
    .A2(\w[35][6] ),
    .A3(\w[39][6] ),
    .S0(net465),
    .S1(net467),
    .X(_03433_));
 sky130_fd_sc_hd__mux4_2 _26703_ (.A0(\w[41][6] ),
    .A1(\w[45][6] ),
    .A2(\w[43][6] ),
    .A3(\w[47][6] ),
    .S0(net465),
    .S1(net467),
    .X(_03434_));
 sky130_fd_sc_hd__mux4_2 _26704_ (.A0(\w[49][6] ),
    .A1(\w[53][6] ),
    .A2(\w[51][6] ),
    .A3(\w[55][6] ),
    .S0(net465),
    .S1(net467),
    .X(_03435_));
 sky130_fd_sc_hd__mux4_2 _26705_ (.A0(\w[57][6] ),
    .A1(\w[61][6] ),
    .A2(\w[59][6] ),
    .A3(\w[63][6] ),
    .S0(net465),
    .S1(net467),
    .X(_03436_));
 sky130_fd_sc_hd__mux4_2 _26706_ (.A0(_03433_),
    .A1(_03434_),
    .A2(_03435_),
    .A3(_03436_),
    .S0(\count16_2[3] ),
    .S1(net543),
    .X(_03437_));
 sky130_fd_sc_hd__mux2i_4 _26707_ (.A0(_03432_),
    .A1(_03437_),
    .S(net453),
    .Y(_11880_));
 sky130_fd_sc_hd__mux4_2 _26708_ (.A0(\w[1][26] ),
    .A1(\w[5][26] ),
    .A2(\w[3][26] ),
    .A3(\w[7][26] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03438_));
 sky130_fd_sc_hd__mux4_2 _26709_ (.A0(\w[9][26] ),
    .A1(\w[13][26] ),
    .A2(\w[11][26] ),
    .A3(\w[15][26] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03439_));
 sky130_fd_sc_hd__mux4_2 _26710_ (.A0(\w[17][26] ),
    .A1(\w[21][26] ),
    .A2(\w[19][26] ),
    .A3(\w[23][26] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03440_));
 sky130_fd_sc_hd__mux4_2 _26711_ (.A0(\w[25][26] ),
    .A1(\w[29][26] ),
    .A2(\w[27][26] ),
    .A3(\w[31][26] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03441_));
 sky130_fd_sc_hd__mux4_2 _26712_ (.A0(_03438_),
    .A1(_03439_),
    .A2(_03440_),
    .A3(_03441_),
    .S0(\count2_2[3] ),
    .S1(net540),
    .X(_03442_));
 sky130_fd_sc_hd__mux4_2 _26713_ (.A0(\w[33][26] ),
    .A1(\w[37][26] ),
    .A2(\w[35][26] ),
    .A3(\w[39][26] ),
    .S0(net424),
    .S1(net429),
    .X(_03443_));
 sky130_fd_sc_hd__mux4_2 _26714_ (.A0(\w[41][26] ),
    .A1(\w[45][26] ),
    .A2(\w[43][26] ),
    .A3(\w[47][26] ),
    .S0(net424),
    .S1(net429),
    .X(_03444_));
 sky130_fd_sc_hd__mux4_2 _26715_ (.A0(\w[49][26] ),
    .A1(\w[53][26] ),
    .A2(\w[51][26] ),
    .A3(\w[55][26] ),
    .S0(net541),
    .S1(net429),
    .X(_03445_));
 sky130_fd_sc_hd__mux4_2 _26716_ (.A0(\w[57][26] ),
    .A1(\w[61][26] ),
    .A2(\w[59][26] ),
    .A3(\w[63][26] ),
    .S0(net424),
    .S1(net429),
    .X(_03446_));
 sky130_fd_sc_hd__mux4_2 _26717_ (.A0(_03443_),
    .A1(_03444_),
    .A2(_03445_),
    .A3(_03446_),
    .S0(net417),
    .S1(net540),
    .X(_03447_));
 sky130_fd_sc_hd__mux2i_4 _26718_ (.A0(_03442_),
    .A1(_03447_),
    .S(net413),
    .Y(_03448_));
 sky130_fd_sc_hd__xnor2_1 _26719_ (.A(_03320_),
    .B(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__xnor2_1 _26720_ (.A(_02788_),
    .B(_03449_),
    .Y(_11885_));
 sky130_fd_sc_hd__mux4_2 _26721_ (.A0(\w[0][14] ),
    .A1(\w[4][14] ),
    .A2(\w[2][14] ),
    .A3(\w[6][14] ),
    .S0(net498),
    .S1(net511),
    .X(_03450_));
 sky130_fd_sc_hd__mux4_2 _26722_ (.A0(\w[8][14] ),
    .A1(\w[12][14] ),
    .A2(\w[10][14] ),
    .A3(\w[14][14] ),
    .S0(net498),
    .S1(net511),
    .X(_03451_));
 sky130_fd_sc_hd__mux4_2 _26723_ (.A0(\w[16][14] ),
    .A1(\w[20][14] ),
    .A2(\w[18][14] ),
    .A3(\w[22][14] ),
    .S0(net498),
    .S1(net511),
    .X(_03452_));
 sky130_fd_sc_hd__mux4_2 _26724_ (.A0(\w[24][14] ),
    .A1(\w[28][14] ),
    .A2(\w[26][14] ),
    .A3(\w[30][14] ),
    .S0(net498),
    .S1(net511),
    .X(_03453_));
 sky130_fd_sc_hd__mux4_2 _26725_ (.A0(_03450_),
    .A1(_03451_),
    .A2(_03452_),
    .A3(_03453_),
    .S0(net496),
    .S1(net494),
    .X(_03454_));
 sky130_fd_sc_hd__mux4_2 _26726_ (.A0(\w[32][14] ),
    .A1(\w[36][14] ),
    .A2(\w[34][14] ),
    .A3(\w[38][14] ),
    .S0(net504),
    .S1(net510),
    .X(_03455_));
 sky130_fd_sc_hd__mux4_2 _26727_ (.A0(\w[40][14] ),
    .A1(\w[44][14] ),
    .A2(\w[42][14] ),
    .A3(\w[46][14] ),
    .S0(net504),
    .S1(net510),
    .X(_03456_));
 sky130_fd_sc_hd__mux4_2 _26728_ (.A0(\w[48][14] ),
    .A1(\w[52][14] ),
    .A2(\w[50][14] ),
    .A3(\w[54][14] ),
    .S0(net504),
    .S1(net510),
    .X(_03457_));
 sky130_fd_sc_hd__mux4_2 _26729_ (.A0(\w[56][14] ),
    .A1(\w[60][14] ),
    .A2(\w[58][14] ),
    .A3(\w[62][14] ),
    .S0(net504),
    .S1(net510),
    .X(_03458_));
 sky130_fd_sc_hd__mux4_2 _26730_ (.A0(_03455_),
    .A1(_03456_),
    .A2(_03457_),
    .A3(_03458_),
    .S0(net548),
    .S1(net494),
    .X(_03459_));
 sky130_fd_sc_hd__mux2i_4 _26731_ (.A0(_03454_),
    .A1(_03459_),
    .S(net492),
    .Y(_03460_));
 sky130_fd_sc_hd__mux4_2 _26732_ (.A0(\w[0][25] ),
    .A1(\w[4][25] ),
    .A2(\w[2][25] ),
    .A3(\w[6][25] ),
    .S0(net503),
    .S1(net509),
    .X(_03461_));
 sky130_fd_sc_hd__mux4_2 _26733_ (.A0(\w[8][25] ),
    .A1(\w[12][25] ),
    .A2(\w[10][25] ),
    .A3(\w[14][25] ),
    .S0(net503),
    .S1(net509),
    .X(_03462_));
 sky130_fd_sc_hd__mux4_2 _26734_ (.A0(\w[16][25] ),
    .A1(\w[20][25] ),
    .A2(\w[18][25] ),
    .A3(\w[22][25] ),
    .S0(net503),
    .S1(net509),
    .X(_03463_));
 sky130_fd_sc_hd__mux4_2 _26735_ (.A0(\w[24][25] ),
    .A1(\w[28][25] ),
    .A2(\w[26][25] ),
    .A3(\w[30][25] ),
    .S0(net503),
    .S1(net509),
    .X(_03464_));
 sky130_fd_sc_hd__mux4_2 _26736_ (.A0(_03461_),
    .A1(_03462_),
    .A2(_03463_),
    .A3(_03464_),
    .S0(net496),
    .S1(net494),
    .X(_03465_));
 sky130_fd_sc_hd__mux4_2 _26737_ (.A0(\w[32][25] ),
    .A1(\w[36][25] ),
    .A2(\w[34][25] ),
    .A3(\w[38][25] ),
    .S0(net502),
    .S1(net508),
    .X(_03466_));
 sky130_fd_sc_hd__mux4_2 _26738_ (.A0(\w[40][25] ),
    .A1(\w[44][25] ),
    .A2(\w[42][25] ),
    .A3(\w[46][25] ),
    .S0(net503),
    .S1(net509),
    .X(_03467_));
 sky130_fd_sc_hd__mux4_2 _26739_ (.A0(\w[48][25] ),
    .A1(\w[52][25] ),
    .A2(\w[50][25] ),
    .A3(\w[54][25] ),
    .S0(net503),
    .S1(net509),
    .X(_03468_));
 sky130_fd_sc_hd__mux4_2 _26740_ (.A0(\w[56][25] ),
    .A1(\w[60][25] ),
    .A2(\w[58][25] ),
    .A3(\w[62][25] ),
    .S0(net503),
    .S1(net509),
    .X(_03469_));
 sky130_fd_sc_hd__mux4_2 _26741_ (.A0(_03466_),
    .A1(_03467_),
    .A2(_03468_),
    .A3(_03469_),
    .S0(net548),
    .S1(net494),
    .X(_03470_));
 sky130_fd_sc_hd__mux2i_4 _26742_ (.A0(_03465_),
    .A1(_03470_),
    .S(net493),
    .Y(_03471_));
 sky130_fd_sc_hd__xnor2_1 _26743_ (.A(_03460_),
    .B(_03471_),
    .Y(_03472_));
 sky130_fd_sc_hd__xnor2_1 _26744_ (.A(_03205_),
    .B(_03472_),
    .Y(_11884_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_53 ();
 sky130_fd_sc_hd__mux4_2 _26746_ (.A0(\w[0][7] ),
    .A1(\w[4][7] ),
    .A2(\w[2][7] ),
    .A3(\w[6][7] ),
    .S0(net380),
    .S1(net388),
    .X(_03474_));
 sky130_fd_sc_hd__mux4_2 _26747_ (.A0(\w[8][7] ),
    .A1(\w[12][7] ),
    .A2(\w[10][7] ),
    .A3(\w[14][7] ),
    .S0(net380),
    .S1(net388),
    .X(_03475_));
 sky130_fd_sc_hd__mux4_2 _26748_ (.A0(\w[16][7] ),
    .A1(\w[20][7] ),
    .A2(\w[18][7] ),
    .A3(\w[22][7] ),
    .S0(net380),
    .S1(net388),
    .X(_03476_));
 sky130_fd_sc_hd__mux4_2 _26749_ (.A0(\w[24][7] ),
    .A1(\w[28][7] ),
    .A2(\w[26][7] ),
    .A3(\w[30][7] ),
    .S0(net380),
    .S1(net388),
    .X(_03477_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_52 ();
 sky130_fd_sc_hd__mux4_2 _26751_ (.A0(_03474_),
    .A1(_03475_),
    .A2(_03476_),
    .A3(_03477_),
    .S0(net379),
    .S1(net376),
    .X(_03479_));
 sky130_fd_sc_hd__mux4_2 _26752_ (.A0(\w[32][7] ),
    .A1(\w[36][7] ),
    .A2(\w[34][7] ),
    .A3(\w[38][7] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_03480_));
 sky130_fd_sc_hd__mux4_2 _26753_ (.A0(\w[40][7] ),
    .A1(\w[44][7] ),
    .A2(\w[42][7] ),
    .A3(\w[46][7] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_03481_));
 sky130_fd_sc_hd__mux4_2 _26754_ (.A0(\w[48][7] ),
    .A1(\w[52][7] ),
    .A2(\w[50][7] ),
    .A3(\w[54][7] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_03482_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_51 ();
 sky130_fd_sc_hd__mux4_2 _26756_ (.A0(\w[56][7] ),
    .A1(\w[60][7] ),
    .A2(\w[58][7] ),
    .A3(\w[62][7] ),
    .S0(\count7_2[2] ),
    .S1(\count7_2[1] ),
    .X(_03484_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_50 ();
 sky130_fd_sc_hd__mux4_2 _26758_ (.A0(_03480_),
    .A1(_03481_),
    .A2(_03482_),
    .A3(_03484_),
    .S0(net379),
    .S1(net376),
    .X(_03486_));
 sky130_fd_sc_hd__mux2i_4 _26759_ (.A0(_03479_),
    .A1(_03486_),
    .S(net373),
    .Y(_11883_));
 sky130_fd_sc_hd__mux4_2 _26760_ (.A0(\w[1][7] ),
    .A1(\w[5][7] ),
    .A2(\w[3][7] ),
    .A3(\w[7][7] ),
    .S0(net461),
    .S1(net544),
    .X(_03487_));
 sky130_fd_sc_hd__mux4_2 _26761_ (.A0(\w[9][7] ),
    .A1(\w[13][7] ),
    .A2(\w[11][7] ),
    .A3(\w[15][7] ),
    .S0(net461),
    .S1(net544),
    .X(_03488_));
 sky130_fd_sc_hd__mux4_2 _26762_ (.A0(\w[17][7] ),
    .A1(\w[21][7] ),
    .A2(\w[19][7] ),
    .A3(\w[23][7] ),
    .S0(net461),
    .S1(net544),
    .X(_03489_));
 sky130_fd_sc_hd__mux4_2 _26763_ (.A0(\w[25][7] ),
    .A1(\w[29][7] ),
    .A2(\w[27][7] ),
    .A3(\w[31][7] ),
    .S0(net461),
    .S1(net544),
    .X(_03490_));
 sky130_fd_sc_hd__mux4_2 _26764_ (.A0(_03487_),
    .A1(_03488_),
    .A2(_03489_),
    .A3(_03490_),
    .S0(net457),
    .S1(\count16_2[4] ),
    .X(_03491_));
 sky130_fd_sc_hd__mux4_2 _26765_ (.A0(\w[33][7] ),
    .A1(\w[37][7] ),
    .A2(\w[35][7] ),
    .A3(\w[39][7] ),
    .S0(net461),
    .S1(net470),
    .X(_03492_));
 sky130_fd_sc_hd__mux4_2 _26766_ (.A0(\w[41][7] ),
    .A1(\w[45][7] ),
    .A2(\w[43][7] ),
    .A3(\w[47][7] ),
    .S0(net461),
    .S1(net470),
    .X(_03493_));
 sky130_fd_sc_hd__mux4_2 _26767_ (.A0(\w[49][7] ),
    .A1(\w[53][7] ),
    .A2(\w[51][7] ),
    .A3(\w[55][7] ),
    .S0(net461),
    .S1(net470),
    .X(_03494_));
 sky130_fd_sc_hd__mux4_2 _26768_ (.A0(\w[57][7] ),
    .A1(\w[61][7] ),
    .A2(\w[59][7] ),
    .A3(\w[63][7] ),
    .S0(net461),
    .S1(net470),
    .X(_03495_));
 sky130_fd_sc_hd__mux4_2 _26769_ (.A0(_03492_),
    .A1(_03493_),
    .A2(_03494_),
    .A3(_03495_),
    .S0(net457),
    .S1(net543),
    .X(_03496_));
 sky130_fd_sc_hd__mux2i_4 _26770_ (.A0(_03491_),
    .A1(_03496_),
    .S(net453),
    .Y(_11888_));
 sky130_fd_sc_hd__mux4_2 _26771_ (.A0(\w[1][27] ),
    .A1(\w[5][27] ),
    .A2(\w[3][27] ),
    .A3(\w[7][27] ),
    .S0(net422),
    .S1(net429),
    .X(_03497_));
 sky130_fd_sc_hd__mux4_2 _26772_ (.A0(\w[9][27] ),
    .A1(\w[13][27] ),
    .A2(\w[11][27] ),
    .A3(\w[15][27] ),
    .S0(net422),
    .S1(net429),
    .X(_03498_));
 sky130_fd_sc_hd__mux4_2 _26773_ (.A0(\w[17][27] ),
    .A1(\w[21][27] ),
    .A2(\w[19][27] ),
    .A3(\w[23][27] ),
    .S0(net422),
    .S1(net429),
    .X(_03499_));
 sky130_fd_sc_hd__mux4_2 _26774_ (.A0(\w[25][27] ),
    .A1(\w[29][27] ),
    .A2(\w[27][27] ),
    .A3(\w[31][27] ),
    .S0(net422),
    .S1(net429),
    .X(_03500_));
 sky130_fd_sc_hd__mux4_2 _26775_ (.A0(_03497_),
    .A1(_03498_),
    .A2(_03499_),
    .A3(_03500_),
    .S0(net416),
    .S1(net414),
    .X(_03501_));
 sky130_fd_sc_hd__mux4_2 _26776_ (.A0(\w[33][27] ),
    .A1(\w[37][27] ),
    .A2(\w[35][27] ),
    .A3(\w[39][27] ),
    .S0(net423),
    .S1(net428),
    .X(_03502_));
 sky130_fd_sc_hd__mux4_2 _26777_ (.A0(\w[41][27] ),
    .A1(\w[45][27] ),
    .A2(\w[43][27] ),
    .A3(\w[47][27] ),
    .S0(net423),
    .S1(net428),
    .X(_03503_));
 sky130_fd_sc_hd__mux4_2 _26778_ (.A0(\w[49][27] ),
    .A1(\w[53][27] ),
    .A2(\w[51][27] ),
    .A3(\w[55][27] ),
    .S0(net423),
    .S1(net428),
    .X(_03504_));
 sky130_fd_sc_hd__mux4_2 _26779_ (.A0(\w[57][27] ),
    .A1(\w[61][27] ),
    .A2(\w[59][27] ),
    .A3(\w[63][27] ),
    .S0(net423),
    .S1(net428),
    .X(_03505_));
 sky130_fd_sc_hd__mux4_2 _26780_ (.A0(_03502_),
    .A1(_03503_),
    .A2(_03504_),
    .A3(_03505_),
    .S0(net417),
    .S1(net414),
    .X(_03506_));
 sky130_fd_sc_hd__mux2i_4 _26781_ (.A0(_03501_),
    .A1(_03506_),
    .S(net413),
    .Y(_03507_));
 sky130_fd_sc_hd__xnor2_1 _26782_ (.A(_03389_),
    .B(_03507_),
    .Y(_03508_));
 sky130_fd_sc_hd__xnor2_1 _26783_ (.A(_02964_),
    .B(_03508_),
    .Y(_11893_));
 sky130_fd_sc_hd__mux4_2 _26784_ (.A0(\w[0][15] ),
    .A1(\w[4][15] ),
    .A2(\w[2][15] ),
    .A3(\w[6][15] ),
    .S0(net1133),
    .S1(net506),
    .X(_03509_));
 sky130_fd_sc_hd__mux4_2 _26785_ (.A0(\w[8][15] ),
    .A1(\w[12][15] ),
    .A2(\w[10][15] ),
    .A3(\w[14][15] ),
    .S0(net1133),
    .S1(net506),
    .X(_03510_));
 sky130_fd_sc_hd__mux4_2 _26786_ (.A0(\w[16][15] ),
    .A1(\w[20][15] ),
    .A2(\w[18][15] ),
    .A3(\w[22][15] ),
    .S0(net1133),
    .S1(net506),
    .X(_03511_));
 sky130_fd_sc_hd__mux4_2 _26787_ (.A0(\w[24][15] ),
    .A1(\w[28][15] ),
    .A2(\w[26][15] ),
    .A3(\w[30][15] ),
    .S0(net1133),
    .S1(net506),
    .X(_03512_));
 sky130_fd_sc_hd__mux4_2 _26788_ (.A0(_03509_),
    .A1(_03510_),
    .A2(_03511_),
    .A3(_03512_),
    .S0(net496),
    .S1(net547),
    .X(_03513_));
 sky130_fd_sc_hd__mux4_2 _26789_ (.A0(\w[32][15] ),
    .A1(\w[36][15] ),
    .A2(\w[34][15] ),
    .A3(\w[38][15] ),
    .S0(net499),
    .S1(net506),
    .X(_03514_));
 sky130_fd_sc_hd__mux4_2 _26790_ (.A0(\w[40][15] ),
    .A1(\w[44][15] ),
    .A2(\w[42][15] ),
    .A3(\w[46][15] ),
    .S0(net499),
    .S1(net506),
    .X(_03515_));
 sky130_fd_sc_hd__mux4_2 _26791_ (.A0(\w[48][15] ),
    .A1(\w[52][15] ),
    .A2(\w[50][15] ),
    .A3(\w[54][15] ),
    .S0(net499),
    .S1(net506),
    .X(_03516_));
 sky130_fd_sc_hd__mux4_2 _26792_ (.A0(\w[56][15] ),
    .A1(\w[60][15] ),
    .A2(\w[58][15] ),
    .A3(\w[62][15] ),
    .S0(net499),
    .S1(net506),
    .X(_03517_));
 sky130_fd_sc_hd__mux4_2 _26793_ (.A0(_03514_),
    .A1(_03515_),
    .A2(_03516_),
    .A3(_03517_),
    .S0(\count15_2[3] ),
    .S1(net547),
    .X(_03518_));
 sky130_fd_sc_hd__mux2i_4 _26794_ (.A0(_03513_),
    .A1(_03518_),
    .S(net493),
    .Y(_03519_));
 sky130_fd_sc_hd__mux4_2 _26795_ (.A0(\w[0][26] ),
    .A1(\w[4][26] ),
    .A2(\w[2][26] ),
    .A3(\w[6][26] ),
    .S0(net498),
    .S1(net509),
    .X(_03520_));
 sky130_fd_sc_hd__mux4_2 _26796_ (.A0(\w[8][26] ),
    .A1(\w[12][26] ),
    .A2(\w[10][26] ),
    .A3(\w[14][26] ),
    .S0(net498),
    .S1(net509),
    .X(_03521_));
 sky130_fd_sc_hd__mux4_2 _26797_ (.A0(\w[16][26] ),
    .A1(\w[20][26] ),
    .A2(\w[18][26] ),
    .A3(\w[22][26] ),
    .S0(net498),
    .S1(net509),
    .X(_03522_));
 sky130_fd_sc_hd__mux4_2 _26798_ (.A0(\w[24][26] ),
    .A1(\w[28][26] ),
    .A2(\w[26][26] ),
    .A3(\w[30][26] ),
    .S0(net498),
    .S1(net509),
    .X(_03523_));
 sky130_fd_sc_hd__mux4_2 _26799_ (.A0(_03520_),
    .A1(_03521_),
    .A2(_03522_),
    .A3(_03523_),
    .S0(net496),
    .S1(net494),
    .X(_03524_));
 sky130_fd_sc_hd__mux4_2 _26800_ (.A0(\w[32][26] ),
    .A1(\w[36][26] ),
    .A2(\w[34][26] ),
    .A3(\w[38][26] ),
    .S0(net503),
    .S1(net509),
    .X(_03525_));
 sky130_fd_sc_hd__mux4_2 _26801_ (.A0(\w[40][26] ),
    .A1(\w[44][26] ),
    .A2(\w[42][26] ),
    .A3(\w[46][26] ),
    .S0(net503),
    .S1(net509),
    .X(_03526_));
 sky130_fd_sc_hd__mux4_2 _26802_ (.A0(\w[48][26] ),
    .A1(\w[52][26] ),
    .A2(\w[50][26] ),
    .A3(\w[54][26] ),
    .S0(net503),
    .S1(net509),
    .X(_03527_));
 sky130_fd_sc_hd__mux4_2 _26803_ (.A0(\w[56][26] ),
    .A1(\w[60][26] ),
    .A2(\w[58][26] ),
    .A3(\w[62][26] ),
    .S0(net503),
    .S1(net509),
    .X(_03528_));
 sky130_fd_sc_hd__mux4_2 _26804_ (.A0(_03525_),
    .A1(_03526_),
    .A2(_03527_),
    .A3(_03528_),
    .S0(net548),
    .S1(net494),
    .X(_03529_));
 sky130_fd_sc_hd__mux2i_4 _26805_ (.A0(_03524_),
    .A1(_03529_),
    .S(net493),
    .Y(_03530_));
 sky130_fd_sc_hd__xnor2_1 _26806_ (.A(_03519_),
    .B(_03530_),
    .Y(_03531_));
 sky130_fd_sc_hd__xnor2_1 _26807_ (.A(_03275_),
    .B(_03531_),
    .Y(_11892_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_49 ();
 sky130_fd_sc_hd__mux4_2 _26809_ (.A0(\w[0][8] ),
    .A1(\w[4][8] ),
    .A2(\w[2][8] ),
    .A3(\w[6][8] ),
    .S0(net382),
    .S1(net389),
    .X(_03533_));
 sky130_fd_sc_hd__mux4_2 _26810_ (.A0(\w[8][8] ),
    .A1(\w[12][8] ),
    .A2(\w[10][8] ),
    .A3(\w[14][8] ),
    .S0(net382),
    .S1(net389),
    .X(_03534_));
 sky130_fd_sc_hd__mux4_2 _26811_ (.A0(\w[16][8] ),
    .A1(\w[20][8] ),
    .A2(\w[18][8] ),
    .A3(\w[22][8] ),
    .S0(net382),
    .S1(net389),
    .X(_03535_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_48 ();
 sky130_fd_sc_hd__mux4_2 _26813_ (.A0(\w[24][8] ),
    .A1(\w[28][8] ),
    .A2(\w[26][8] ),
    .A3(\w[30][8] ),
    .S0(net382),
    .S1(net389),
    .X(_03537_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_47 ();
 sky130_fd_sc_hd__mux4_2 _26815_ (.A0(_03533_),
    .A1(_03534_),
    .A2(_03535_),
    .A3(_03537_),
    .S0(net377),
    .S1(net375),
    .X(_03539_));
 sky130_fd_sc_hd__mux4_2 _26816_ (.A0(\w[32][8] ),
    .A1(\w[36][8] ),
    .A2(\w[34][8] ),
    .A3(\w[38][8] ),
    .S0(net382),
    .S1(net389),
    .X(_03540_));
 sky130_fd_sc_hd__mux4_2 _26817_ (.A0(\w[40][8] ),
    .A1(\w[44][8] ),
    .A2(\w[42][8] ),
    .A3(\w[46][8] ),
    .S0(net382),
    .S1(net389),
    .X(_03541_));
 sky130_fd_sc_hd__mux4_2 _26818_ (.A0(\w[48][8] ),
    .A1(\w[52][8] ),
    .A2(\w[50][8] ),
    .A3(\w[54][8] ),
    .S0(net382),
    .S1(net389),
    .X(_03542_));
 sky130_fd_sc_hd__mux4_2 _26819_ (.A0(\w[56][8] ),
    .A1(\w[60][8] ),
    .A2(\w[58][8] ),
    .A3(\w[62][8] ),
    .S0(net383),
    .S1(net390),
    .X(_03543_));
 sky130_fd_sc_hd__mux4_2 _26820_ (.A0(_03540_),
    .A1(_03541_),
    .A2(_03542_),
    .A3(_03543_),
    .S0(net378),
    .S1(net535),
    .X(_03544_));
 sky130_fd_sc_hd__mux2i_4 _26821_ (.A0(_03539_),
    .A1(_03544_),
    .S(net374),
    .Y(_11891_));
 sky130_fd_sc_hd__mux4_2 _26822_ (.A0(\w[1][8] ),
    .A1(\w[5][8] ),
    .A2(\w[3][8] ),
    .A3(\w[7][8] ),
    .S0(net464),
    .S1(net468),
    .X(_03545_));
 sky130_fd_sc_hd__mux4_2 _26823_ (.A0(\w[9][8] ),
    .A1(\w[13][8] ),
    .A2(\w[11][8] ),
    .A3(\w[15][8] ),
    .S0(net464),
    .S1(net468),
    .X(_03546_));
 sky130_fd_sc_hd__mux4_2 _26824_ (.A0(\w[17][8] ),
    .A1(\w[21][8] ),
    .A2(\w[19][8] ),
    .A3(\w[23][8] ),
    .S0(net464),
    .S1(net468),
    .X(_03547_));
 sky130_fd_sc_hd__mux4_2 _26825_ (.A0(\w[25][8] ),
    .A1(\w[29][8] ),
    .A2(\w[27][8] ),
    .A3(\w[31][8] ),
    .S0(net464),
    .S1(net468),
    .X(_03548_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_46 ();
 sky130_fd_sc_hd__mux4_2 _26827_ (.A0(_03545_),
    .A1(_03546_),
    .A2(_03547_),
    .A3(_03548_),
    .S0(\count16_2[3] ),
    .S1(net454),
    .X(_03550_));
 sky130_fd_sc_hd__mux4_2 _26828_ (.A0(\w[33][8] ),
    .A1(\w[37][8] ),
    .A2(\w[35][8] ),
    .A3(\w[39][8] ),
    .S0(net464),
    .S1(net467),
    .X(_03551_));
 sky130_fd_sc_hd__mux4_2 _26829_ (.A0(\w[41][8] ),
    .A1(\w[45][8] ),
    .A2(\w[43][8] ),
    .A3(\w[47][8] ),
    .S0(net464),
    .S1(net467),
    .X(_03552_));
 sky130_fd_sc_hd__mux4_2 _26830_ (.A0(\w[49][8] ),
    .A1(\w[53][8] ),
    .A2(\w[51][8] ),
    .A3(\w[55][8] ),
    .S0(net464),
    .S1(net467),
    .X(_03553_));
 sky130_fd_sc_hd__mux4_2 _26831_ (.A0(\w[57][8] ),
    .A1(\w[61][8] ),
    .A2(\w[59][8] ),
    .A3(\w[63][8] ),
    .S0(net464),
    .S1(net467),
    .X(_03554_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_45 ();
 sky130_fd_sc_hd__mux4_2 _26833_ (.A0(_03551_),
    .A1(_03552_),
    .A2(_03553_),
    .A3(_03554_),
    .S0(\count16_2[3] ),
    .S1(net543),
    .X(_03556_));
 sky130_fd_sc_hd__mux2i_4 _26834_ (.A0(_03550_),
    .A1(_03556_),
    .S(net542),
    .Y(_11896_));
 sky130_fd_sc_hd__mux4_2 _26835_ (.A0(\w[1][28] ),
    .A1(\w[5][28] ),
    .A2(\w[3][28] ),
    .A3(\w[7][28] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03557_));
 sky130_fd_sc_hd__mux4_2 _26836_ (.A0(\w[9][28] ),
    .A1(\w[13][28] ),
    .A2(\w[11][28] ),
    .A3(\w[15][28] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03558_));
 sky130_fd_sc_hd__mux4_2 _26837_ (.A0(\w[17][28] ),
    .A1(\w[21][28] ),
    .A2(\w[19][28] ),
    .A3(\w[23][28] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03559_));
 sky130_fd_sc_hd__mux4_2 _26838_ (.A0(\w[25][28] ),
    .A1(\w[29][28] ),
    .A2(\w[27][28] ),
    .A3(\w[31][28] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03560_));
 sky130_fd_sc_hd__mux4_2 _26839_ (.A0(_03557_),
    .A1(_03558_),
    .A2(_03559_),
    .A3(_03560_),
    .S0(\count2_2[3] ),
    .S1(net540),
    .X(_03561_));
 sky130_fd_sc_hd__mux4_2 _26840_ (.A0(\w[33][28] ),
    .A1(\w[37][28] ),
    .A2(\w[35][28] ),
    .A3(\w[39][28] ),
    .S0(net541),
    .S1(net431),
    .X(_03562_));
 sky130_fd_sc_hd__mux4_2 _26841_ (.A0(\w[41][28] ),
    .A1(\w[45][28] ),
    .A2(\w[43][28] ),
    .A3(\w[47][28] ),
    .S0(net541),
    .S1(net431),
    .X(_03563_));
 sky130_fd_sc_hd__mux4_2 _26842_ (.A0(\w[49][28] ),
    .A1(\w[53][28] ),
    .A2(\w[51][28] ),
    .A3(\w[55][28] ),
    .S0(net541),
    .S1(net431),
    .X(_03564_));
 sky130_fd_sc_hd__mux4_2 _26843_ (.A0(\w[57][28] ),
    .A1(\w[61][28] ),
    .A2(\w[59][28] ),
    .A3(\w[63][28] ),
    .S0(net541),
    .S1(net431),
    .X(_03565_));
 sky130_fd_sc_hd__mux4_2 _26844_ (.A0(_03562_),
    .A1(_03563_),
    .A2(_03564_),
    .A3(_03565_),
    .S0(\count2_2[3] ),
    .S1(net540),
    .X(_03566_));
 sky130_fd_sc_hd__mux2i_4 _26845_ (.A0(_03561_),
    .A1(_03566_),
    .S(net413),
    .Y(_03567_));
 sky130_fd_sc_hd__xnor2_1 _26846_ (.A(_03448_),
    .B(_03567_),
    .Y(_03568_));
 sky130_fd_sc_hd__xnor2_1 _26847_ (.A(_02770_),
    .B(_03568_),
    .Y(_11901_));
 sky130_fd_sc_hd__mux4_2 _26848_ (.A0(\w[0][16] ),
    .A1(\w[4][16] ),
    .A2(\w[2][16] ),
    .A3(\w[6][16] ),
    .S0(net1133),
    .S1(net506),
    .X(_03569_));
 sky130_fd_sc_hd__mux4_2 _26849_ (.A0(\w[8][16] ),
    .A1(\w[12][16] ),
    .A2(\w[10][16] ),
    .A3(\w[14][16] ),
    .S0(net1133),
    .S1(\count15_2[1] ),
    .X(_03570_));
 sky130_fd_sc_hd__mux4_2 _26850_ (.A0(\w[16][16] ),
    .A1(\w[20][16] ),
    .A2(\w[18][16] ),
    .A3(\w[22][16] ),
    .S0(net1133),
    .S1(\count15_2[1] ),
    .X(_03571_));
 sky130_fd_sc_hd__mux4_2 _26851_ (.A0(\w[24][16] ),
    .A1(\w[28][16] ),
    .A2(\w[26][16] ),
    .A3(\w[30][16] ),
    .S0(net1133),
    .S1(\count15_2[1] ),
    .X(_03572_));
 sky130_fd_sc_hd__mux4_2 _26852_ (.A0(_03569_),
    .A1(_03570_),
    .A2(_03571_),
    .A3(_03572_),
    .S0(\count15_2[3] ),
    .S1(\count15_2[4] ),
    .X(_03573_));
 sky130_fd_sc_hd__mux4_2 _26853_ (.A0(\w[32][16] ),
    .A1(\w[36][16] ),
    .A2(\w[34][16] ),
    .A3(\w[38][16] ),
    .S0(net505),
    .S1(net511),
    .X(_03574_));
 sky130_fd_sc_hd__mux4_2 _26854_ (.A0(\w[40][16] ),
    .A1(\w[44][16] ),
    .A2(\w[42][16] ),
    .A3(\w[46][16] ),
    .S0(net505),
    .S1(net511),
    .X(_03575_));
 sky130_fd_sc_hd__mux4_2 _26855_ (.A0(\w[48][16] ),
    .A1(\w[52][16] ),
    .A2(\w[50][16] ),
    .A3(\w[54][16] ),
    .S0(net505),
    .S1(net511),
    .X(_03576_));
 sky130_fd_sc_hd__mux4_2 _26856_ (.A0(\w[56][16] ),
    .A1(\w[60][16] ),
    .A2(\w[58][16] ),
    .A3(\w[62][16] ),
    .S0(net505),
    .S1(net511),
    .X(_03577_));
 sky130_fd_sc_hd__mux4_2 _26857_ (.A0(_03574_),
    .A1(_03575_),
    .A2(_03576_),
    .A3(_03577_),
    .S0(net497),
    .S1(net495),
    .X(_03578_));
 sky130_fd_sc_hd__mux2i_4 _26858_ (.A0(_03573_),
    .A1(_03578_),
    .S(\count15_2[5] ),
    .Y(_03579_));
 sky130_fd_sc_hd__mux4_2 _26859_ (.A0(\w[0][27] ),
    .A1(\w[4][27] ),
    .A2(\w[2][27] ),
    .A3(\w[6][27] ),
    .S0(net498),
    .S1(net511),
    .X(_03580_));
 sky130_fd_sc_hd__mux4_2 _26860_ (.A0(\w[8][27] ),
    .A1(\w[12][27] ),
    .A2(\w[10][27] ),
    .A3(\w[14][27] ),
    .S0(net498),
    .S1(net511),
    .X(_03581_));
 sky130_fd_sc_hd__mux4_2 _26861_ (.A0(\w[16][27] ),
    .A1(\w[20][27] ),
    .A2(\w[18][27] ),
    .A3(\w[22][27] ),
    .S0(net498),
    .S1(net511),
    .X(_03582_));
 sky130_fd_sc_hd__mux4_2 _26862_ (.A0(\w[24][27] ),
    .A1(\w[28][27] ),
    .A2(\w[26][27] ),
    .A3(\w[30][27] ),
    .S0(net498),
    .S1(net511),
    .X(_03583_));
 sky130_fd_sc_hd__mux4_2 _26863_ (.A0(_03580_),
    .A1(_03581_),
    .A2(_03582_),
    .A3(_03583_),
    .S0(net496),
    .S1(net494),
    .X(_03584_));
 sky130_fd_sc_hd__mux4_2 _26864_ (.A0(\w[32][27] ),
    .A1(\w[36][27] ),
    .A2(\w[34][27] ),
    .A3(\w[38][27] ),
    .S0(net499),
    .S1(net511),
    .X(_03585_));
 sky130_fd_sc_hd__mux4_2 _26865_ (.A0(\w[40][27] ),
    .A1(\w[44][27] ),
    .A2(\w[42][27] ),
    .A3(\w[46][27] ),
    .S0(net499),
    .S1(net511),
    .X(_03586_));
 sky130_fd_sc_hd__mux4_2 _26866_ (.A0(\w[48][27] ),
    .A1(\w[52][27] ),
    .A2(\w[50][27] ),
    .A3(\w[54][27] ),
    .S0(net499),
    .S1(net511),
    .X(_03587_));
 sky130_fd_sc_hd__mux4_2 _26867_ (.A0(\w[56][27] ),
    .A1(\w[60][27] ),
    .A2(\w[58][27] ),
    .A3(\w[62][27] ),
    .S0(net499),
    .S1(net511),
    .X(_03588_));
 sky130_fd_sc_hd__mux4_2 _26868_ (.A0(_03585_),
    .A1(_03586_),
    .A2(_03587_),
    .A3(_03588_),
    .S0(net496),
    .S1(net547),
    .X(_03589_));
 sky130_fd_sc_hd__mux2i_4 _26869_ (.A0(_03584_),
    .A1(_03589_),
    .S(net493),
    .Y(_03590_));
 sky130_fd_sc_hd__xnor2_1 _26870_ (.A(_03579_),
    .B(_03590_),
    .Y(_03591_));
 sky130_fd_sc_hd__xnor2_1 _26871_ (.A(_03344_),
    .B(_03591_),
    .Y(_11900_));
 sky130_fd_sc_hd__mux4_2 _26872_ (.A0(\w[0][9] ),
    .A1(\w[4][9] ),
    .A2(\w[2][9] ),
    .A3(\w[6][9] ),
    .S0(net381),
    .S1(net389),
    .X(_03592_));
 sky130_fd_sc_hd__mux4_2 _26873_ (.A0(\w[8][9] ),
    .A1(\w[12][9] ),
    .A2(\w[10][9] ),
    .A3(\w[14][9] ),
    .S0(net381),
    .S1(net389),
    .X(_03593_));
 sky130_fd_sc_hd__mux4_2 _26874_ (.A0(\w[16][9] ),
    .A1(\w[20][9] ),
    .A2(\w[18][9] ),
    .A3(\w[22][9] ),
    .S0(net381),
    .S1(net389),
    .X(_03594_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_44 ();
 sky130_fd_sc_hd__mux4_2 _26876_ (.A0(\w[24][9] ),
    .A1(\w[28][9] ),
    .A2(\w[26][9] ),
    .A3(\w[30][9] ),
    .S0(net381),
    .S1(net389),
    .X(_03596_));
 sky130_fd_sc_hd__mux4_2 _26877_ (.A0(_03592_),
    .A1(_03593_),
    .A2(_03594_),
    .A3(_03596_),
    .S0(net378),
    .S1(net535),
    .X(_03597_));
 sky130_fd_sc_hd__mux4_2 _26878_ (.A0(\w[32][9] ),
    .A1(\w[36][9] ),
    .A2(\w[34][9] ),
    .A3(\w[38][9] ),
    .S0(net383),
    .S1(net390),
    .X(_03598_));
 sky130_fd_sc_hd__mux4_2 _26879_ (.A0(\w[40][9] ),
    .A1(\w[44][9] ),
    .A2(\w[42][9] ),
    .A3(\w[46][9] ),
    .S0(net383),
    .S1(net390),
    .X(_03599_));
 sky130_fd_sc_hd__mux4_2 _26880_ (.A0(\w[48][9] ),
    .A1(\w[52][9] ),
    .A2(\w[50][9] ),
    .A3(\w[54][9] ),
    .S0(net383),
    .S1(net390),
    .X(_03600_));
 sky130_fd_sc_hd__mux4_2 _26881_ (.A0(\w[56][9] ),
    .A1(\w[60][9] ),
    .A2(\w[58][9] ),
    .A3(\w[62][9] ),
    .S0(net383),
    .S1(net390),
    .X(_03601_));
 sky130_fd_sc_hd__mux4_2 _26882_ (.A0(_03598_),
    .A1(_03599_),
    .A2(_03600_),
    .A3(_03601_),
    .S0(net378),
    .S1(net535),
    .X(_03602_));
 sky130_fd_sc_hd__mux2i_4 _26883_ (.A0(_03597_),
    .A1(_03602_),
    .S(net374),
    .Y(_11899_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_43 ();
 sky130_fd_sc_hd__mux4_2 _26885_ (.A0(\w[1][9] ),
    .A1(\w[5][9] ),
    .A2(\w[3][9] ),
    .A3(\w[7][9] ),
    .S0(net462),
    .S1(net471),
    .X(_03604_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_42 ();
 sky130_fd_sc_hd__mux4_2 _26887_ (.A0(\w[9][9] ),
    .A1(\w[13][9] ),
    .A2(\w[11][9] ),
    .A3(\w[15][9] ),
    .S0(net462),
    .S1(net471),
    .X(_03606_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_41 ();
 sky130_fd_sc_hd__mux4_2 _26889_ (.A0(\w[17][9] ),
    .A1(\w[21][9] ),
    .A2(\w[19][9] ),
    .A3(\w[23][9] ),
    .S0(net462),
    .S1(net471),
    .X(_03608_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_40 ();
 sky130_fd_sc_hd__mux4_2 _26891_ (.A0(\w[25][9] ),
    .A1(\w[29][9] ),
    .A2(\w[27][9] ),
    .A3(\w[31][9] ),
    .S0(net462),
    .S1(net471),
    .X(_03610_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_39 ();
 sky130_fd_sc_hd__mux4_2 _26893_ (.A0(_03604_),
    .A1(_03606_),
    .A2(_03608_),
    .A3(_03610_),
    .S0(net457),
    .S1(\count16_2[4] ),
    .X(_03612_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_38 ();
 sky130_fd_sc_hd__mux4_2 _26895_ (.A0(\w[33][9] ),
    .A1(\w[37][9] ),
    .A2(\w[35][9] ),
    .A3(\w[39][9] ),
    .S0(net461),
    .S1(net471),
    .X(_03614_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_37 ();
 sky130_fd_sc_hd__mux4_2 _26897_ (.A0(\w[41][9] ),
    .A1(\w[45][9] ),
    .A2(\w[43][9] ),
    .A3(\w[47][9] ),
    .S0(net461),
    .S1(net471),
    .X(_03616_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_36 ();
 sky130_fd_sc_hd__mux4_2 _26899_ (.A0(\w[49][9] ),
    .A1(\w[53][9] ),
    .A2(\w[51][9] ),
    .A3(\w[55][9] ),
    .S0(net461),
    .S1(net471),
    .X(_03618_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_35 ();
 sky130_fd_sc_hd__mux4_2 _26901_ (.A0(\w[57][9] ),
    .A1(\w[61][9] ),
    .A2(\w[59][9] ),
    .A3(\w[63][9] ),
    .S0(net461),
    .S1(net471),
    .X(_03620_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_34 ();
 sky130_fd_sc_hd__mux4_2 _26903_ (.A0(_03614_),
    .A1(_03616_),
    .A2(_03618_),
    .A3(_03620_),
    .S0(net457),
    .S1(net543),
    .X(_03622_));
 sky130_fd_sc_hd__mux2i_4 _26904_ (.A0(_03612_),
    .A1(_03622_),
    .S(net542),
    .Y(_11904_));
 sky130_fd_sc_hd__mux4_2 _26905_ (.A0(\w[1][29] ),
    .A1(\w[5][29] ),
    .A2(\w[3][29] ),
    .A3(\w[7][29] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03623_));
 sky130_fd_sc_hd__mux4_2 _26906_ (.A0(\w[9][29] ),
    .A1(\w[13][29] ),
    .A2(\w[11][29] ),
    .A3(\w[15][29] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03624_));
 sky130_fd_sc_hd__mux4_2 _26907_ (.A0(\w[17][29] ),
    .A1(\w[21][29] ),
    .A2(\w[19][29] ),
    .A3(\w[23][29] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03625_));
 sky130_fd_sc_hd__mux4_2 _26908_ (.A0(\w[25][29] ),
    .A1(\w[29][29] ),
    .A2(\w[27][29] ),
    .A3(\w[31][29] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03626_));
 sky130_fd_sc_hd__mux4_2 _26909_ (.A0(_03623_),
    .A1(_03624_),
    .A2(_03625_),
    .A3(_03626_),
    .S0(\count2_2[3] ),
    .S1(net540),
    .X(_03627_));
 sky130_fd_sc_hd__mux4_2 _26910_ (.A0(\w[33][29] ),
    .A1(\w[37][29] ),
    .A2(\w[35][29] ),
    .A3(\w[39][29] ),
    .S0(net425),
    .S1(net430),
    .X(_03628_));
 sky130_fd_sc_hd__mux4_2 _26911_ (.A0(\w[41][29] ),
    .A1(\w[45][29] ),
    .A2(\w[43][29] ),
    .A3(\w[47][29] ),
    .S0(net425),
    .S1(net430),
    .X(_03629_));
 sky130_fd_sc_hd__mux4_2 _26912_ (.A0(\w[49][29] ),
    .A1(\w[53][29] ),
    .A2(\w[51][29] ),
    .A3(\w[55][29] ),
    .S0(net425),
    .S1(net430),
    .X(_03630_));
 sky130_fd_sc_hd__mux4_2 _26913_ (.A0(\w[57][29] ),
    .A1(\w[61][29] ),
    .A2(\w[59][29] ),
    .A3(\w[63][29] ),
    .S0(net425),
    .S1(net430),
    .X(_03631_));
 sky130_fd_sc_hd__mux4_2 _26914_ (.A0(_03628_),
    .A1(_03629_),
    .A2(_03630_),
    .A3(_03631_),
    .S0(net417),
    .S1(net540),
    .X(_03632_));
 sky130_fd_sc_hd__mux2i_4 _26915_ (.A0(_03627_),
    .A1(_03632_),
    .S(\count2_2[5] ),
    .Y(_03633_));
 sky130_fd_sc_hd__xnor2_1 _26916_ (.A(_03507_),
    .B(_03633_),
    .Y(_03634_));
 sky130_fd_sc_hd__xnor2_1 _26917_ (.A(_02953_),
    .B(_03634_),
    .Y(_11909_));
 sky130_fd_sc_hd__mux4_2 _26918_ (.A0(\w[0][28] ),
    .A1(\w[4][28] ),
    .A2(\w[2][28] ),
    .A3(\w[6][28] ),
    .S0(net498),
    .S1(net511),
    .X(_03635_));
 sky130_fd_sc_hd__mux4_2 _26919_ (.A0(\w[8][28] ),
    .A1(\w[12][28] ),
    .A2(\w[10][28] ),
    .A3(\w[14][28] ),
    .S0(net498),
    .S1(net511),
    .X(_03636_));
 sky130_fd_sc_hd__mux4_2 _26920_ (.A0(\w[16][28] ),
    .A1(\w[20][28] ),
    .A2(\w[18][28] ),
    .A3(\w[22][28] ),
    .S0(net498),
    .S1(net511),
    .X(_03637_));
 sky130_fd_sc_hd__mux4_2 _26921_ (.A0(\w[24][28] ),
    .A1(\w[28][28] ),
    .A2(\w[26][28] ),
    .A3(\w[30][28] ),
    .S0(net498),
    .S1(net511),
    .X(_03638_));
 sky130_fd_sc_hd__mux4_2 _26922_ (.A0(_03635_),
    .A1(_03636_),
    .A2(_03637_),
    .A3(_03638_),
    .S0(net496),
    .S1(net494),
    .X(_03639_));
 sky130_fd_sc_hd__mux4_2 _26923_ (.A0(\w[32][28] ),
    .A1(\w[36][28] ),
    .A2(\w[34][28] ),
    .A3(\w[38][28] ),
    .S0(net503),
    .S1(net509),
    .X(_03640_));
 sky130_fd_sc_hd__mux4_2 _26924_ (.A0(\w[40][28] ),
    .A1(\w[44][28] ),
    .A2(\w[42][28] ),
    .A3(\w[46][28] ),
    .S0(net503),
    .S1(net509),
    .X(_03641_));
 sky130_fd_sc_hd__mux4_2 _26925_ (.A0(\w[48][28] ),
    .A1(\w[52][28] ),
    .A2(\w[50][28] ),
    .A3(\w[54][28] ),
    .S0(net503),
    .S1(net509),
    .X(_03642_));
 sky130_fd_sc_hd__mux4_2 _26926_ (.A0(\w[56][28] ),
    .A1(\w[60][28] ),
    .A2(\w[58][28] ),
    .A3(\w[62][28] ),
    .S0(net503),
    .S1(net509),
    .X(_03643_));
 sky130_fd_sc_hd__mux4_2 _26927_ (.A0(_03640_),
    .A1(_03641_),
    .A2(_03642_),
    .A3(_03643_),
    .S0(\count15_2[3] ),
    .S1(net494),
    .X(_03644_));
 sky130_fd_sc_hd__mux2i_4 _26928_ (.A0(_03639_),
    .A1(_03644_),
    .S(net493),
    .Y(_03645_));
 sky130_fd_sc_hd__mux4_2 _26929_ (.A0(\w[0][17] ),
    .A1(\w[4][17] ),
    .A2(\w[2][17] ),
    .A3(\w[6][17] ),
    .S0(net498),
    .S1(net511),
    .X(_03646_));
 sky130_fd_sc_hd__mux4_2 _26930_ (.A0(\w[8][17] ),
    .A1(\w[12][17] ),
    .A2(\w[10][17] ),
    .A3(\w[14][17] ),
    .S0(net498),
    .S1(net511),
    .X(_03647_));
 sky130_fd_sc_hd__mux4_2 _26931_ (.A0(\w[16][17] ),
    .A1(\w[20][17] ),
    .A2(\w[18][17] ),
    .A3(\w[22][17] ),
    .S0(net498),
    .S1(net511),
    .X(_03648_));
 sky130_fd_sc_hd__mux4_2 _26932_ (.A0(\w[24][17] ),
    .A1(\w[28][17] ),
    .A2(\w[26][17] ),
    .A3(\w[30][17] ),
    .S0(net498),
    .S1(net511),
    .X(_03649_));
 sky130_fd_sc_hd__mux4_2 _26933_ (.A0(_03646_),
    .A1(_03647_),
    .A2(_03648_),
    .A3(_03649_),
    .S0(net496),
    .S1(net494),
    .X(_03650_));
 sky130_fd_sc_hd__mux4_2 _26934_ (.A0(\w[32][17] ),
    .A1(\w[36][17] ),
    .A2(\w[34][17] ),
    .A3(\w[38][17] ),
    .S0(net503),
    .S1(net509),
    .X(_03651_));
 sky130_fd_sc_hd__mux4_2 _26935_ (.A0(\w[40][17] ),
    .A1(\w[44][17] ),
    .A2(\w[42][17] ),
    .A3(\w[46][17] ),
    .S0(net503),
    .S1(net509),
    .X(_03652_));
 sky130_fd_sc_hd__mux4_2 _26936_ (.A0(\w[48][17] ),
    .A1(\w[52][17] ),
    .A2(\w[50][17] ),
    .A3(\w[54][17] ),
    .S0(net503),
    .S1(net509),
    .X(_03653_));
 sky130_fd_sc_hd__mux4_2 _26937_ (.A0(\w[56][17] ),
    .A1(\w[60][17] ),
    .A2(\w[58][17] ),
    .A3(\w[62][17] ),
    .S0(net503),
    .S1(net509),
    .X(_03654_));
 sky130_fd_sc_hd__mux4_2 _26938_ (.A0(_03651_),
    .A1(_03652_),
    .A2(_03653_),
    .A3(_03654_),
    .S0(net548),
    .S1(net494),
    .X(_03655_));
 sky130_fd_sc_hd__mux2i_4 _26939_ (.A0(_03650_),
    .A1(_03655_),
    .S(net493),
    .Y(_03656_));
 sky130_fd_sc_hd__xnor2_1 _26940_ (.A(_03645_),
    .B(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__xnor2_1 _26941_ (.A(_03402_),
    .B(_03657_),
    .Y(_11908_));
 sky130_fd_sc_hd__mux4_2 _26942_ (.A0(\w[0][10] ),
    .A1(\w[4][10] ),
    .A2(\w[2][10] ),
    .A3(\w[6][10] ),
    .S0(net381),
    .S1(net389),
    .X(_03658_));
 sky130_fd_sc_hd__mux4_2 _26943_ (.A0(\w[8][10] ),
    .A1(\w[12][10] ),
    .A2(\w[10][10] ),
    .A3(\w[14][10] ),
    .S0(net381),
    .S1(net389),
    .X(_03659_));
 sky130_fd_sc_hd__mux4_2 _26944_ (.A0(\w[16][10] ),
    .A1(\w[20][10] ),
    .A2(\w[18][10] ),
    .A3(\w[22][10] ),
    .S0(net381),
    .S1(net389),
    .X(_03660_));
 sky130_fd_sc_hd__mux4_2 _26945_ (.A0(\w[24][10] ),
    .A1(\w[28][10] ),
    .A2(\w[26][10] ),
    .A3(\w[30][10] ),
    .S0(net381),
    .S1(net389),
    .X(_03661_));
 sky130_fd_sc_hd__mux4_2 _26946_ (.A0(_03658_),
    .A1(_03659_),
    .A2(_03660_),
    .A3(_03661_),
    .S0(net378),
    .S1(net535),
    .X(_03662_));
 sky130_fd_sc_hd__mux4_2 _26947_ (.A0(\w[32][10] ),
    .A1(\w[36][10] ),
    .A2(\w[34][10] ),
    .A3(\w[38][10] ),
    .S0(net383),
    .S1(net390),
    .X(_03663_));
 sky130_fd_sc_hd__mux4_2 _26948_ (.A0(\w[40][10] ),
    .A1(\w[44][10] ),
    .A2(\w[42][10] ),
    .A3(\w[46][10] ),
    .S0(net383),
    .S1(net390),
    .X(_03664_));
 sky130_fd_sc_hd__mux4_2 _26949_ (.A0(\w[48][10] ),
    .A1(\w[52][10] ),
    .A2(\w[50][10] ),
    .A3(\w[54][10] ),
    .S0(net383),
    .S1(net390),
    .X(_03665_));
 sky130_fd_sc_hd__mux4_2 _26950_ (.A0(\w[56][10] ),
    .A1(\w[60][10] ),
    .A2(\w[58][10] ),
    .A3(\w[62][10] ),
    .S0(net383),
    .S1(net390),
    .X(_03666_));
 sky130_fd_sc_hd__mux4_2 _26951_ (.A0(_03663_),
    .A1(_03664_),
    .A2(_03665_),
    .A3(_03666_),
    .S0(net378),
    .S1(net535),
    .X(_03667_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_33 ();
 sky130_fd_sc_hd__mux2i_4 _26953_ (.A0(_03662_),
    .A1(_03667_),
    .S(net374),
    .Y(_11907_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_32 ();
 sky130_fd_sc_hd__mux4_2 _26955_ (.A0(\w[1][10] ),
    .A1(\w[5][10] ),
    .A2(\w[3][10] ),
    .A3(\w[7][10] ),
    .S0(net463),
    .S1(net467),
    .X(_03670_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_31 ();
 sky130_fd_sc_hd__mux4_2 _26957_ (.A0(\w[9][10] ),
    .A1(\w[13][10] ),
    .A2(\w[11][10] ),
    .A3(\w[15][10] ),
    .S0(net463),
    .S1(net467),
    .X(_03672_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_30 ();
 sky130_fd_sc_hd__mux4_2 _26959_ (.A0(\w[17][10] ),
    .A1(\w[21][10] ),
    .A2(\w[19][10] ),
    .A3(\w[23][10] ),
    .S0(net463),
    .S1(net467),
    .X(_03674_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_29 ();
 sky130_fd_sc_hd__mux4_2 _26961_ (.A0(\w[25][10] ),
    .A1(\w[29][10] ),
    .A2(\w[27][10] ),
    .A3(\w[31][10] ),
    .S0(net463),
    .S1(net467),
    .X(_03676_));
 sky130_fd_sc_hd__mux4_2 _26962_ (.A0(_03670_),
    .A1(_03672_),
    .A2(_03674_),
    .A3(_03676_),
    .S0(net458),
    .S1(net455),
    .X(_03677_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_28 ();
 sky130_fd_sc_hd__mux4_2 _26964_ (.A0(\w[33][10] ),
    .A1(\w[37][10] ),
    .A2(\w[35][10] ),
    .A3(\w[39][10] ),
    .S0(net465),
    .S1(net469),
    .X(_03679_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_27 ();
 sky130_fd_sc_hd__mux4_2 _26966_ (.A0(\w[41][10] ),
    .A1(\w[45][10] ),
    .A2(\w[43][10] ),
    .A3(\w[47][10] ),
    .S0(net465),
    .S1(net469),
    .X(_03681_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_26 ();
 sky130_fd_sc_hd__mux4_2 _26968_ (.A0(\w[49][10] ),
    .A1(\w[53][10] ),
    .A2(\w[51][10] ),
    .A3(\w[55][10] ),
    .S0(net464),
    .S1(net469),
    .X(_03683_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_25 ();
 sky130_fd_sc_hd__mux4_2 _26970_ (.A0(\w[57][10] ),
    .A1(\w[61][10] ),
    .A2(\w[59][10] ),
    .A3(\w[63][10] ),
    .S0(net465),
    .S1(net469),
    .X(_03685_));
 sky130_fd_sc_hd__mux4_2 _26971_ (.A0(_03679_),
    .A1(_03681_),
    .A2(_03683_),
    .A3(_03685_),
    .S0(net458),
    .S1(net455),
    .X(_03686_));
 sky130_fd_sc_hd__mux2i_4 _26972_ (.A0(_03677_),
    .A1(_03686_),
    .S(net542),
    .Y(_11912_));
 sky130_fd_sc_hd__mux4_2 _26973_ (.A0(\w[1][30] ),
    .A1(\w[5][30] ),
    .A2(\w[3][30] ),
    .A3(\w[7][30] ),
    .S0(net541),
    .S1(net431),
    .X(_03687_));
 sky130_fd_sc_hd__mux4_2 _26974_ (.A0(\w[9][30] ),
    .A1(\w[13][30] ),
    .A2(\w[11][30] ),
    .A3(\w[15][30] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03688_));
 sky130_fd_sc_hd__mux4_2 _26975_ (.A0(\w[17][30] ),
    .A1(\w[21][30] ),
    .A2(\w[19][30] ),
    .A3(\w[23][30] ),
    .S0(net541),
    .S1(\count2_2[1] ),
    .X(_03689_));
 sky130_fd_sc_hd__mux4_2 _26976_ (.A0(\w[25][30] ),
    .A1(\w[29][30] ),
    .A2(\w[27][30] ),
    .A3(\w[31][30] ),
    .S0(net541),
    .S1(net431),
    .X(_03690_));
 sky130_fd_sc_hd__mux4_2 _26977_ (.A0(_03687_),
    .A1(_03688_),
    .A2(_03689_),
    .A3(_03690_),
    .S0(\count2_2[3] ),
    .S1(\count2_2[4] ),
    .X(_03691_));
 sky130_fd_sc_hd__mux4_2 _26978_ (.A0(\w[33][30] ),
    .A1(\w[37][30] ),
    .A2(\w[35][30] ),
    .A3(\w[39][30] ),
    .S0(net425),
    .S1(net430),
    .X(_03692_));
 sky130_fd_sc_hd__mux4_2 _26979_ (.A0(\w[41][30] ),
    .A1(\w[45][30] ),
    .A2(\w[43][30] ),
    .A3(\w[47][30] ),
    .S0(net425),
    .S1(net430),
    .X(_03693_));
 sky130_fd_sc_hd__mux4_2 _26980_ (.A0(\w[49][30] ),
    .A1(\w[53][30] ),
    .A2(\w[51][30] ),
    .A3(\w[55][30] ),
    .S0(net425),
    .S1(net430),
    .X(_03694_));
 sky130_fd_sc_hd__mux4_2 _26981_ (.A0(\w[57][30] ),
    .A1(\w[61][30] ),
    .A2(\w[59][30] ),
    .A3(\w[63][30] ),
    .S0(net425),
    .S1(net430),
    .X(_03695_));
 sky130_fd_sc_hd__mux4_2 _26982_ (.A0(_03692_),
    .A1(_03693_),
    .A2(_03694_),
    .A3(_03695_),
    .S0(net418),
    .S1(net415),
    .X(_03696_));
 sky130_fd_sc_hd__mux2i_4 _26983_ (.A0(_03691_),
    .A1(_03696_),
    .S(\count2_2[5] ),
    .Y(_03697_));
 sky130_fd_sc_hd__xnor2_1 _26984_ (.A(_03567_),
    .B(_03697_),
    .Y(_03698_));
 sky130_fd_sc_hd__xnor2_2 _26985_ (.A(_03086_),
    .B(_03698_),
    .Y(_11917_));
 sky130_fd_sc_hd__mux4_2 _26986_ (.A0(\w[0][29] ),
    .A1(\w[4][29] ),
    .A2(\w[2][29] ),
    .A3(\w[6][29] ),
    .S0(net498),
    .S1(net506),
    .X(_03699_));
 sky130_fd_sc_hd__mux4_2 _26987_ (.A0(\w[8][29] ),
    .A1(\w[12][29] ),
    .A2(\w[10][29] ),
    .A3(\w[14][29] ),
    .S0(net498),
    .S1(net506),
    .X(_03700_));
 sky130_fd_sc_hd__mux4_2 _26988_ (.A0(\w[16][29] ),
    .A1(\w[20][29] ),
    .A2(\w[18][29] ),
    .A3(\w[22][29] ),
    .S0(net498),
    .S1(net506),
    .X(_03701_));
 sky130_fd_sc_hd__mux4_2 _26989_ (.A0(\w[24][29] ),
    .A1(\w[28][29] ),
    .A2(\w[26][29] ),
    .A3(\w[30][29] ),
    .S0(net498),
    .S1(net506),
    .X(_03702_));
 sky130_fd_sc_hd__mux4_2 _26990_ (.A0(_03699_),
    .A1(_03700_),
    .A2(_03701_),
    .A3(_03702_),
    .S0(net496),
    .S1(net547),
    .X(_03703_));
 sky130_fd_sc_hd__mux4_2 _26991_ (.A0(\w[32][29] ),
    .A1(\w[36][29] ),
    .A2(\w[34][29] ),
    .A3(\w[38][29] ),
    .S0(net499),
    .S1(net506),
    .X(_03704_));
 sky130_fd_sc_hd__mux4_2 _26992_ (.A0(\w[40][29] ),
    .A1(\w[44][29] ),
    .A2(\w[42][29] ),
    .A3(\w[46][29] ),
    .S0(net499),
    .S1(net506),
    .X(_03705_));
 sky130_fd_sc_hd__mux4_2 _26993_ (.A0(\w[48][29] ),
    .A1(\w[52][29] ),
    .A2(\w[50][29] ),
    .A3(\w[54][29] ),
    .S0(net499),
    .S1(net506),
    .X(_03706_));
 sky130_fd_sc_hd__mux4_2 _26994_ (.A0(\w[56][29] ),
    .A1(\w[60][29] ),
    .A2(\w[58][29] ),
    .A3(\w[62][29] ),
    .S0(net499),
    .S1(net506),
    .X(_03707_));
 sky130_fd_sc_hd__mux4_2 _26995_ (.A0(_03704_),
    .A1(_03705_),
    .A2(_03706_),
    .A3(_03707_),
    .S0(net496),
    .S1(net547),
    .X(_03708_));
 sky130_fd_sc_hd__mux2i_4 _26996_ (.A0(_03703_),
    .A1(_03708_),
    .S(net493),
    .Y(_03709_));
 sky130_fd_sc_hd__xnor2_1 _26997_ (.A(_03460_),
    .B(_03709_),
    .Y(_03710_));
 sky130_fd_sc_hd__xnor2_1 _26998_ (.A(_02853_),
    .B(_03710_),
    .Y(_11916_));
 sky130_fd_sc_hd__mux4_2 _26999_ (.A0(\w[0][11] ),
    .A1(\w[4][11] ),
    .A2(\w[2][11] ),
    .A3(\w[6][11] ),
    .S0(net382),
    .S1(net389),
    .X(_03711_));
 sky130_fd_sc_hd__mux4_2 _27000_ (.A0(\w[8][11] ),
    .A1(\w[12][11] ),
    .A2(\w[10][11] ),
    .A3(\w[14][11] ),
    .S0(net382),
    .S1(net389),
    .X(_03712_));
 sky130_fd_sc_hd__mux4_2 _27001_ (.A0(\w[16][11] ),
    .A1(\w[20][11] ),
    .A2(\w[18][11] ),
    .A3(\w[22][11] ),
    .S0(net382),
    .S1(net389),
    .X(_03713_));
 sky130_fd_sc_hd__mux4_2 _27002_ (.A0(\w[24][11] ),
    .A1(\w[28][11] ),
    .A2(\w[26][11] ),
    .A3(\w[30][11] ),
    .S0(net382),
    .S1(net389),
    .X(_03714_));
 sky130_fd_sc_hd__mux4_2 _27003_ (.A0(_03711_),
    .A1(_03712_),
    .A2(_03713_),
    .A3(_03714_),
    .S0(net377),
    .S1(net375),
    .X(_03715_));
 sky130_fd_sc_hd__mux4_2 _27004_ (.A0(\w[32][11] ),
    .A1(\w[36][11] ),
    .A2(\w[34][11] ),
    .A3(\w[38][11] ),
    .S0(net385),
    .S1(net392),
    .X(_03716_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_24 ();
 sky130_fd_sc_hd__mux4_2 _27006_ (.A0(\w[40][11] ),
    .A1(\w[44][11] ),
    .A2(\w[42][11] ),
    .A3(\w[46][11] ),
    .S0(net385),
    .S1(net392),
    .X(_03718_));
 sky130_fd_sc_hd__mux4_2 _27007_ (.A0(\w[48][11] ),
    .A1(\w[52][11] ),
    .A2(\w[50][11] ),
    .A3(\w[54][11] ),
    .S0(net385),
    .S1(net392),
    .X(_03719_));
 sky130_fd_sc_hd__mux4_2 _27008_ (.A0(\w[56][11] ),
    .A1(\w[60][11] ),
    .A2(\w[58][11] ),
    .A3(\w[62][11] ),
    .S0(net385),
    .S1(net392),
    .X(_03720_));
 sky130_fd_sc_hd__mux4_2 _27009_ (.A0(_03716_),
    .A1(_03718_),
    .A2(_03719_),
    .A3(_03720_),
    .S0(net378),
    .S1(\count7_2[4] ),
    .X(_03721_));
 sky130_fd_sc_hd__mux2i_2 _27010_ (.A0(_03715_),
    .A1(_03721_),
    .S(net374),
    .Y(_11915_));
 sky130_fd_sc_hd__mux4_2 _27011_ (.A0(\w[1][11] ),
    .A1(\w[5][11] ),
    .A2(\w[3][11] ),
    .A3(\w[7][11] ),
    .S0(net464),
    .S1(net468),
    .X(_03722_));
 sky130_fd_sc_hd__mux4_2 _27012_ (.A0(\w[9][11] ),
    .A1(\w[13][11] ),
    .A2(\w[11][11] ),
    .A3(\w[15][11] ),
    .S0(net464),
    .S1(net468),
    .X(_03723_));
 sky130_fd_sc_hd__mux4_2 _27013_ (.A0(\w[17][11] ),
    .A1(\w[21][11] ),
    .A2(\w[19][11] ),
    .A3(\w[23][11] ),
    .S0(net464),
    .S1(net468),
    .X(_03724_));
 sky130_fd_sc_hd__mux4_2 _27014_ (.A0(\w[25][11] ),
    .A1(\w[29][11] ),
    .A2(\w[27][11] ),
    .A3(\w[31][11] ),
    .S0(net464),
    .S1(net468),
    .X(_03725_));
 sky130_fd_sc_hd__mux4_2 _27015_ (.A0(_03722_),
    .A1(_03723_),
    .A2(_03724_),
    .A3(_03725_),
    .S0(\count16_2[3] ),
    .S1(net454),
    .X(_03726_));
 sky130_fd_sc_hd__mux4_2 _27016_ (.A0(\w[33][11] ),
    .A1(\w[37][11] ),
    .A2(\w[35][11] ),
    .A3(\w[39][11] ),
    .S0(\count16_2[2] ),
    .S1(net471),
    .X(_03727_));
 sky130_fd_sc_hd__mux4_2 _27017_ (.A0(\w[41][11] ),
    .A1(\w[45][11] ),
    .A2(\w[43][11] ),
    .A3(\w[47][11] ),
    .S0(\count16_2[2] ),
    .S1(net471),
    .X(_03728_));
 sky130_fd_sc_hd__mux4_2 _27018_ (.A0(\w[49][11] ),
    .A1(\w[53][11] ),
    .A2(\w[51][11] ),
    .A3(\w[55][11] ),
    .S0(\count16_2[2] ),
    .S1(net471),
    .X(_03729_));
 sky130_fd_sc_hd__mux4_2 _27019_ (.A0(\w[57][11] ),
    .A1(\w[61][11] ),
    .A2(\w[59][11] ),
    .A3(\w[63][11] ),
    .S0(\count16_2[2] ),
    .S1(net471),
    .X(_03730_));
 sky130_fd_sc_hd__mux4_2 _27020_ (.A0(_03727_),
    .A1(_03728_),
    .A2(_03729_),
    .A3(_03730_),
    .S0(net458),
    .S1(net455),
    .X(_03731_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_23 ();
 sky130_fd_sc_hd__mux2i_2 _27022_ (.A0(_03726_),
    .A1(_03731_),
    .S(net542),
    .Y(_11920_));
 sky130_fd_sc_hd__mux4_2 _27023_ (.A0(\w[1][31] ),
    .A1(\w[5][31] ),
    .A2(\w[3][31] ),
    .A3(\w[7][31] ),
    .S0(net422),
    .S1(net431),
    .X(_03733_));
 sky130_fd_sc_hd__mux4_2 _27024_ (.A0(\w[9][31] ),
    .A1(\w[13][31] ),
    .A2(\w[11][31] ),
    .A3(\w[15][31] ),
    .S0(net422),
    .S1(net431),
    .X(_03734_));
 sky130_fd_sc_hd__mux4_2 _27025_ (.A0(\w[17][31] ),
    .A1(\w[21][31] ),
    .A2(\w[19][31] ),
    .A3(\w[23][31] ),
    .S0(net422),
    .S1(net431),
    .X(_03735_));
 sky130_fd_sc_hd__mux4_2 _27026_ (.A0(\w[25][31] ),
    .A1(\w[29][31] ),
    .A2(\w[27][31] ),
    .A3(\w[31][31] ),
    .S0(net422),
    .S1(net431),
    .X(_03736_));
 sky130_fd_sc_hd__mux4_2 _27027_ (.A0(_03733_),
    .A1(_03734_),
    .A2(_03735_),
    .A3(_03736_),
    .S0(net417),
    .S1(net414),
    .X(_03737_));
 sky130_fd_sc_hd__mux4_2 _27028_ (.A0(\w[33][31] ),
    .A1(\w[37][31] ),
    .A2(\w[35][31] ),
    .A3(\w[39][31] ),
    .S0(net424),
    .S1(net429),
    .X(_03738_));
 sky130_fd_sc_hd__mux4_2 _27029_ (.A0(\w[41][31] ),
    .A1(\w[45][31] ),
    .A2(\w[43][31] ),
    .A3(\w[47][31] ),
    .S0(net424),
    .S1(net429),
    .X(_03739_));
 sky130_fd_sc_hd__mux4_2 _27030_ (.A0(\w[49][31] ),
    .A1(\w[53][31] ),
    .A2(\w[51][31] ),
    .A3(\w[55][31] ),
    .S0(net424),
    .S1(net429),
    .X(_03740_));
 sky130_fd_sc_hd__mux4_2 _27031_ (.A0(\w[57][31] ),
    .A1(\w[61][31] ),
    .A2(\w[59][31] ),
    .A3(\w[63][31] ),
    .S0(net424),
    .S1(net429),
    .X(_03741_));
 sky130_fd_sc_hd__mux4_2 _27032_ (.A0(_03738_),
    .A1(_03739_),
    .A2(_03740_),
    .A3(_03741_),
    .S0(net417),
    .S1(net540),
    .X(_03742_));
 sky130_fd_sc_hd__mux2i_4 _27033_ (.A0(_03737_),
    .A1(_03742_),
    .S(net413),
    .Y(_03743_));
 sky130_fd_sc_hd__xnor2_1 _27034_ (.A(_03633_),
    .B(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__xnor2_1 _27035_ (.A(_03168_),
    .B(_03744_),
    .Y(_11925_));
 sky130_fd_sc_hd__mux4_2 _27036_ (.A0(\w[0][30] ),
    .A1(\w[4][30] ),
    .A2(\w[2][30] ),
    .A3(\w[6][30] ),
    .S0(net499),
    .S1(net506),
    .X(_03745_));
 sky130_fd_sc_hd__mux4_2 _27037_ (.A0(\w[8][30] ),
    .A1(\w[12][30] ),
    .A2(\w[10][30] ),
    .A3(\w[14][30] ),
    .S0(net499),
    .S1(net506),
    .X(_03746_));
 sky130_fd_sc_hd__mux4_2 _27038_ (.A0(\w[16][30] ),
    .A1(\w[20][30] ),
    .A2(\w[18][30] ),
    .A3(\w[22][30] ),
    .S0(net499),
    .S1(net506),
    .X(_03747_));
 sky130_fd_sc_hd__mux4_2 _27039_ (.A0(\w[24][30] ),
    .A1(\w[28][30] ),
    .A2(\w[26][30] ),
    .A3(\w[30][30] ),
    .S0(net499),
    .S1(net506),
    .X(_03748_));
 sky130_fd_sc_hd__mux4_2 _27040_ (.A0(_03745_),
    .A1(_03746_),
    .A2(_03747_),
    .A3(_03748_),
    .S0(net496),
    .S1(net547),
    .X(_03749_));
 sky130_fd_sc_hd__mux4_2 _27041_ (.A0(\w[32][30] ),
    .A1(\w[36][30] ),
    .A2(\w[34][30] ),
    .A3(\w[38][30] ),
    .S0(net499),
    .S1(net506),
    .X(_03750_));
 sky130_fd_sc_hd__mux4_2 _27042_ (.A0(\w[40][30] ),
    .A1(\w[44][30] ),
    .A2(\w[42][30] ),
    .A3(\w[46][30] ),
    .S0(net499),
    .S1(net506),
    .X(_03751_));
 sky130_fd_sc_hd__mux4_2 _27043_ (.A0(\w[48][30] ),
    .A1(\w[52][30] ),
    .A2(\w[50][30] ),
    .A3(\w[54][30] ),
    .S0(net499),
    .S1(net506),
    .X(_03752_));
 sky130_fd_sc_hd__mux4_2 _27044_ (.A0(\w[56][30] ),
    .A1(\w[60][30] ),
    .A2(\w[58][30] ),
    .A3(\w[62][30] ),
    .S0(net499),
    .S1(net506),
    .X(_03753_));
 sky130_fd_sc_hd__mux4_2 _27045_ (.A0(_03750_),
    .A1(_03751_),
    .A2(_03752_),
    .A3(_03753_),
    .S0(net496),
    .S1(net547),
    .X(_03754_));
 sky130_fd_sc_hd__mux2i_4 _27046_ (.A0(_03749_),
    .A1(_03754_),
    .S(net493),
    .Y(_03755_));
 sky130_fd_sc_hd__xnor2_1 _27047_ (.A(_03519_),
    .B(_03755_),
    .Y(_03756_));
 sky130_fd_sc_hd__xnor2_1 _27048_ (.A(_03005_),
    .B(_03756_),
    .Y(_11924_));
 sky130_fd_sc_hd__mux4_2 _27049_ (.A0(\w[0][12] ),
    .A1(\w[4][12] ),
    .A2(\w[2][12] ),
    .A3(\w[6][12] ),
    .S0(net386),
    .S1(net393),
    .X(_03757_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_22 ();
 sky130_fd_sc_hd__mux4_2 _27051_ (.A0(\w[8][12] ),
    .A1(\w[12][12] ),
    .A2(\w[10][12] ),
    .A3(\w[14][12] ),
    .S0(net386),
    .S1(net393),
    .X(_03759_));
 sky130_fd_sc_hd__mux4_2 _27052_ (.A0(\w[16][12] ),
    .A1(\w[20][12] ),
    .A2(\w[18][12] ),
    .A3(\w[22][12] ),
    .S0(net386),
    .S1(net393),
    .X(_03760_));
 sky130_fd_sc_hd__mux4_2 _27053_ (.A0(\w[24][12] ),
    .A1(\w[28][12] ),
    .A2(\w[26][12] ),
    .A3(\w[30][12] ),
    .S0(net386),
    .S1(net393),
    .X(_03761_));
 sky130_fd_sc_hd__mux4_2 _27054_ (.A0(_03757_),
    .A1(_03759_),
    .A2(_03760_),
    .A3(_03761_),
    .S0(net379),
    .S1(net376),
    .X(_03762_));
 sky130_fd_sc_hd__mux4_2 _27055_ (.A0(\w[32][12] ),
    .A1(\w[36][12] ),
    .A2(\w[34][12] ),
    .A3(\w[38][12] ),
    .S0(net386),
    .S1(net393),
    .X(_03763_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_21 ();
 sky130_fd_sc_hd__mux4_2 _27057_ (.A0(\w[40][12] ),
    .A1(\w[44][12] ),
    .A2(\w[42][12] ),
    .A3(\w[46][12] ),
    .S0(net386),
    .S1(net393),
    .X(_03765_));
 sky130_fd_sc_hd__mux4_2 _27058_ (.A0(\w[48][12] ),
    .A1(\w[52][12] ),
    .A2(\w[50][12] ),
    .A3(\w[54][12] ),
    .S0(net386),
    .S1(net393),
    .X(_03766_));
 sky130_fd_sc_hd__mux4_2 _27059_ (.A0(\w[56][12] ),
    .A1(\w[60][12] ),
    .A2(\w[58][12] ),
    .A3(\w[62][12] ),
    .S0(net386),
    .S1(net393),
    .X(_03767_));
 sky130_fd_sc_hd__mux4_2 _27060_ (.A0(_03763_),
    .A1(_03765_),
    .A2(_03766_),
    .A3(_03767_),
    .S0(net379),
    .S1(net376),
    .X(_03768_));
 sky130_fd_sc_hd__mux2i_4 _27061_ (.A0(_03762_),
    .A1(_03768_),
    .S(net373),
    .Y(_11923_));
 sky130_fd_sc_hd__mux4_2 _27062_ (.A0(\w[1][12] ),
    .A1(\w[5][12] ),
    .A2(\w[3][12] ),
    .A3(\w[7][12] ),
    .S0(net465),
    .S1(net468),
    .X(_03769_));
 sky130_fd_sc_hd__mux4_2 _27063_ (.A0(\w[9][12] ),
    .A1(\w[13][12] ),
    .A2(\w[11][12] ),
    .A3(\w[15][12] ),
    .S0(net465),
    .S1(net468),
    .X(_03770_));
 sky130_fd_sc_hd__mux4_2 _27064_ (.A0(\w[17][12] ),
    .A1(\w[21][12] ),
    .A2(\w[19][12] ),
    .A3(\w[23][12] ),
    .S0(net465),
    .S1(net468),
    .X(_03771_));
 sky130_fd_sc_hd__mux4_2 _27065_ (.A0(\w[25][12] ),
    .A1(\w[29][12] ),
    .A2(\w[27][12] ),
    .A3(\w[31][12] ),
    .S0(net465),
    .S1(net468),
    .X(_03772_));
 sky130_fd_sc_hd__mux4_2 _27066_ (.A0(_03769_),
    .A1(_03770_),
    .A2(_03771_),
    .A3(_03772_),
    .S0(net458),
    .S1(net455),
    .X(_03773_));
 sky130_fd_sc_hd__mux4_2 _27067_ (.A0(\w[33][12] ),
    .A1(\w[37][12] ),
    .A2(\w[35][12] ),
    .A3(\w[39][12] ),
    .S0(net465),
    .S1(net469),
    .X(_03774_));
 sky130_fd_sc_hd__mux4_2 _27068_ (.A0(\w[41][12] ),
    .A1(\w[45][12] ),
    .A2(\w[43][12] ),
    .A3(\w[47][12] ),
    .S0(net465),
    .S1(net469),
    .X(_03775_));
 sky130_fd_sc_hd__mux4_2 _27069_ (.A0(\w[49][12] ),
    .A1(\w[53][12] ),
    .A2(\w[51][12] ),
    .A3(\w[55][12] ),
    .S0(net465),
    .S1(net469),
    .X(_03776_));
 sky130_fd_sc_hd__mux4_2 _27070_ (.A0(\w[57][12] ),
    .A1(\w[61][12] ),
    .A2(\w[59][12] ),
    .A3(\w[63][12] ),
    .S0(net465),
    .S1(net469),
    .X(_03777_));
 sky130_fd_sc_hd__mux4_2 _27071_ (.A0(_03774_),
    .A1(_03775_),
    .A2(_03776_),
    .A3(_03777_),
    .S0(net458),
    .S1(net455),
    .X(_03778_));
 sky130_fd_sc_hd__mux2i_4 _27072_ (.A0(_03773_),
    .A1(_03778_),
    .S(net542),
    .Y(_11928_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_19 ();
 sky130_fd_sc_hd__mux4_2 _27075_ (.A0(\w[1][0] ),
    .A1(\w[5][0] ),
    .A2(\w[3][0] ),
    .A3(\w[7][0] ),
    .S0(net422),
    .S1(net429),
    .X(_03781_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_17 ();
 sky130_fd_sc_hd__mux4_2 _27078_ (.A0(\w[9][0] ),
    .A1(\w[13][0] ),
    .A2(\w[11][0] ),
    .A3(\w[15][0] ),
    .S0(net422),
    .S1(net429),
    .X(_03784_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_15 ();
 sky130_fd_sc_hd__mux4_2 _27081_ (.A0(\w[17][0] ),
    .A1(\w[21][0] ),
    .A2(\w[19][0] ),
    .A3(\w[23][0] ),
    .S0(net422),
    .S1(net429),
    .X(_03787_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_13 ();
 sky130_fd_sc_hd__mux4_2 _27084_ (.A0(\w[25][0] ),
    .A1(\w[29][0] ),
    .A2(\w[27][0] ),
    .A3(\w[31][0] ),
    .S0(net422),
    .S1(net429),
    .X(_03790_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_11 ();
 sky130_fd_sc_hd__mux4_2 _27087_ (.A0(_03781_),
    .A1(_03784_),
    .A2(_03787_),
    .A3(_03790_),
    .S0(net416),
    .S1(net414),
    .X(_03793_));
 sky130_fd_sc_hd__mux4_2 _27088_ (.A0(\w[33][0] ),
    .A1(\w[37][0] ),
    .A2(\w[35][0] ),
    .A3(\w[39][0] ),
    .S0(net423),
    .S1(net428),
    .X(_03794_));
 sky130_fd_sc_hd__mux4_2 _27089_ (.A0(\w[41][0] ),
    .A1(\w[45][0] ),
    .A2(\w[43][0] ),
    .A3(\w[47][0] ),
    .S0(net423),
    .S1(net428),
    .X(_03795_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_9 ();
 sky130_fd_sc_hd__mux4_2 _27092_ (.A0(\w[49][0] ),
    .A1(\w[53][0] ),
    .A2(\w[51][0] ),
    .A3(\w[55][0] ),
    .S0(net423),
    .S1(net428),
    .X(_03798_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_7 ();
 sky130_fd_sc_hd__mux4_2 _27095_ (.A0(\w[57][0] ),
    .A1(\w[61][0] ),
    .A2(\w[59][0] ),
    .A3(\w[63][0] ),
    .S0(net423),
    .S1(net428),
    .X(_03801_));
 sky130_fd_sc_hd__mux4_2 _27096_ (.A0(_03794_),
    .A1(_03795_),
    .A2(_03798_),
    .A3(_03801_),
    .S0(net416),
    .S1(net414),
    .X(_03802_));
 sky130_fd_sc_hd__mux2i_4 _27097_ (.A0(_03793_),
    .A1(_03802_),
    .S(net413),
    .Y(_03803_));
 sky130_fd_sc_hd__xnor2_1 _27098_ (.A(_03697_),
    .B(_03803_),
    .Y(_03804_));
 sky130_fd_sc_hd__xnor2_1 _27099_ (.A(_03250_),
    .B(_03804_),
    .Y(_11933_));
 sky130_fd_sc_hd__mux4_2 _27100_ (.A0(\w[0][31] ),
    .A1(\w[4][31] ),
    .A2(\w[2][31] ),
    .A3(\w[6][31] ),
    .S0(net503),
    .S1(net509),
    .X(_03805_));
 sky130_fd_sc_hd__mux4_2 _27101_ (.A0(\w[8][31] ),
    .A1(\w[12][31] ),
    .A2(\w[10][31] ),
    .A3(\w[14][31] ),
    .S0(net503),
    .S1(net509),
    .X(_03806_));
 sky130_fd_sc_hd__mux4_2 _27102_ (.A0(\w[16][31] ),
    .A1(\w[20][31] ),
    .A2(\w[18][31] ),
    .A3(\w[22][31] ),
    .S0(net503),
    .S1(net509),
    .X(_03807_));
 sky130_fd_sc_hd__mux4_2 _27103_ (.A0(\w[24][31] ),
    .A1(\w[28][31] ),
    .A2(\w[26][31] ),
    .A3(\w[30][31] ),
    .S0(net503),
    .S1(net509),
    .X(_03808_));
 sky130_fd_sc_hd__mux4_2 _27104_ (.A0(_03805_),
    .A1(_03806_),
    .A2(_03807_),
    .A3(_03808_),
    .S0(net496),
    .S1(net494),
    .X(_03809_));
 sky130_fd_sc_hd__mux4_2 _27105_ (.A0(\w[32][31] ),
    .A1(\w[36][31] ),
    .A2(\w[34][31] ),
    .A3(\w[38][31] ),
    .S0(net502),
    .S1(net508),
    .X(_03810_));
 sky130_fd_sc_hd__mux4_2 _27106_ (.A0(\w[40][31] ),
    .A1(\w[44][31] ),
    .A2(\w[42][31] ),
    .A3(\w[46][31] ),
    .S0(net502),
    .S1(net508),
    .X(_03811_));
 sky130_fd_sc_hd__mux4_2 _27107_ (.A0(\w[48][31] ),
    .A1(\w[52][31] ),
    .A2(\w[50][31] ),
    .A3(\w[54][31] ),
    .S0(net502),
    .S1(net508),
    .X(_03812_));
 sky130_fd_sc_hd__mux4_2 _27108_ (.A0(\w[56][31] ),
    .A1(\w[60][31] ),
    .A2(\w[58][31] ),
    .A3(\w[62][31] ),
    .S0(net504),
    .S1(net510),
    .X(_03813_));
 sky130_fd_sc_hd__mux4_2 _27109_ (.A0(_03810_),
    .A1(_03811_),
    .A2(_03812_),
    .A3(_03813_),
    .S0(net548),
    .S1(net494),
    .X(_03814_));
 sky130_fd_sc_hd__mux2i_4 _27110_ (.A0(_03809_),
    .A1(_03814_),
    .S(net492),
    .Y(_03815_));
 sky130_fd_sc_hd__xnor2_1 _27111_ (.A(_03579_),
    .B(_03815_),
    .Y(_03816_));
 sky130_fd_sc_hd__xnor2_1 _27112_ (.A(_03109_),
    .B(_03816_),
    .Y(_11932_));
 sky130_fd_sc_hd__mux4_2 _27113_ (.A0(\w[0][13] ),
    .A1(\w[4][13] ),
    .A2(\w[2][13] ),
    .A3(\w[6][13] ),
    .S0(net384),
    .S1(net391),
    .X(_03817_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_6 ();
 sky130_fd_sc_hd__mux4_2 _27115_ (.A0(\w[8][13] ),
    .A1(\w[12][13] ),
    .A2(\w[10][13] ),
    .A3(\w[14][13] ),
    .S0(net384),
    .S1(net391),
    .X(_03819_));
 sky130_fd_sc_hd__mux4_2 _27116_ (.A0(\w[16][13] ),
    .A1(\w[20][13] ),
    .A2(\w[18][13] ),
    .A3(\w[22][13] ),
    .S0(net384),
    .S1(net391),
    .X(_03820_));
 sky130_fd_sc_hd__mux4_2 _27117_ (.A0(\w[24][13] ),
    .A1(\w[28][13] ),
    .A2(\w[26][13] ),
    .A3(\w[30][13] ),
    .S0(net384),
    .S1(net391),
    .X(_03821_));
 sky130_fd_sc_hd__mux4_2 _27118_ (.A0(_03817_),
    .A1(_03819_),
    .A2(_03820_),
    .A3(_03821_),
    .S0(net377),
    .S1(net375),
    .X(_03822_));
 sky130_fd_sc_hd__mux4_2 _27119_ (.A0(\w[32][13] ),
    .A1(\w[36][13] ),
    .A2(\w[34][13] ),
    .A3(\w[38][13] ),
    .S0(net385),
    .S1(net392),
    .X(_03823_));
 sky130_fd_sc_hd__mux4_2 _27120_ (.A0(\w[40][13] ),
    .A1(\w[44][13] ),
    .A2(\w[42][13] ),
    .A3(\w[46][13] ),
    .S0(net385),
    .S1(net392),
    .X(_03824_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_5 ();
 sky130_fd_sc_hd__mux4_2 _27122_ (.A0(\w[48][13] ),
    .A1(\w[52][13] ),
    .A2(\w[50][13] ),
    .A3(\w[54][13] ),
    .S0(net386),
    .S1(net393),
    .X(_03826_));
 sky130_fd_sc_hd__mux4_2 _27123_ (.A0(\w[56][13] ),
    .A1(\w[60][13] ),
    .A2(\w[58][13] ),
    .A3(\w[62][13] ),
    .S0(\count7_2[2] ),
    .S1(net393),
    .X(_03827_));
 sky130_fd_sc_hd__mux4_2 _27124_ (.A0(_03823_),
    .A1(_03824_),
    .A2(_03826_),
    .A3(_03827_),
    .S0(net379),
    .S1(net376),
    .X(_03828_));
 sky130_fd_sc_hd__mux2i_4 _27125_ (.A0(_03822_),
    .A1(_03828_),
    .S(net373),
    .Y(_11931_));
 sky130_fd_sc_hd__mux4_2 _27126_ (.A0(\w[1][13] ),
    .A1(\w[5][13] ),
    .A2(\w[3][13] ),
    .A3(\w[7][13] ),
    .S0(net463),
    .S1(net467),
    .X(_03829_));
 sky130_fd_sc_hd__mux4_2 _27127_ (.A0(\w[9][13] ),
    .A1(\w[13][13] ),
    .A2(\w[11][13] ),
    .A3(\w[15][13] ),
    .S0(net463),
    .S1(net467),
    .X(_03830_));
 sky130_fd_sc_hd__mux4_2 _27128_ (.A0(\w[17][13] ),
    .A1(\w[21][13] ),
    .A2(\w[19][13] ),
    .A3(\w[23][13] ),
    .S0(net463),
    .S1(net467),
    .X(_03831_));
 sky130_fd_sc_hd__mux4_2 _27129_ (.A0(\w[25][13] ),
    .A1(\w[29][13] ),
    .A2(\w[27][13] ),
    .A3(\w[31][13] ),
    .S0(net463),
    .S1(net467),
    .X(_03832_));
 sky130_fd_sc_hd__mux4_2 _27130_ (.A0(_03829_),
    .A1(_03830_),
    .A2(_03831_),
    .A3(_03832_),
    .S0(net458),
    .S1(net455),
    .X(_03833_));
 sky130_fd_sc_hd__mux4_2 _27131_ (.A0(\w[33][13] ),
    .A1(\w[37][13] ),
    .A2(\w[35][13] ),
    .A3(\w[39][13] ),
    .S0(\count16_2[2] ),
    .S1(net471),
    .X(_03834_));
 sky130_fd_sc_hd__mux4_2 _27132_ (.A0(\w[41][13] ),
    .A1(\w[45][13] ),
    .A2(\w[43][13] ),
    .A3(\w[47][13] ),
    .S0(\count16_2[2] ),
    .S1(net471),
    .X(_03835_));
 sky130_fd_sc_hd__mux4_2 _27133_ (.A0(\w[49][13] ),
    .A1(\w[53][13] ),
    .A2(\w[51][13] ),
    .A3(\w[55][13] ),
    .S0(\count16_2[2] ),
    .S1(net471),
    .X(_03836_));
 sky130_fd_sc_hd__mux4_2 _27134_ (.A0(\w[57][13] ),
    .A1(\w[61][13] ),
    .A2(\w[59][13] ),
    .A3(\w[63][13] ),
    .S0(\count16_2[2] ),
    .S1(net471),
    .X(_03837_));
 sky130_fd_sc_hd__mux4_2 _27135_ (.A0(_03834_),
    .A1(_03835_),
    .A2(_03836_),
    .A3(_03837_),
    .S0(net458),
    .S1(net455),
    .X(_03838_));
 sky130_fd_sc_hd__mux2i_4 _27136_ (.A0(_03833_),
    .A1(_03838_),
    .S(net542),
    .Y(_11936_));
 sky130_fd_sc_hd__mux4_2 _27137_ (.A0(\w[1][1] ),
    .A1(\w[5][1] ),
    .A2(\w[3][1] ),
    .A3(\w[7][1] ),
    .S0(net422),
    .S1(net429),
    .X(_03839_));
 sky130_fd_sc_hd__mux4_2 _27138_ (.A0(\w[9][1] ),
    .A1(\w[13][1] ),
    .A2(\w[11][1] ),
    .A3(\w[15][1] ),
    .S0(net422),
    .S1(net431),
    .X(_03840_));
 sky130_fd_sc_hd__mux4_2 _27139_ (.A0(\w[17][1] ),
    .A1(\w[21][1] ),
    .A2(\w[19][1] ),
    .A3(\w[23][1] ),
    .S0(net422),
    .S1(net429),
    .X(_03841_));
 sky130_fd_sc_hd__mux4_2 _27140_ (.A0(\w[25][1] ),
    .A1(\w[29][1] ),
    .A2(\w[27][1] ),
    .A3(\w[31][1] ),
    .S0(net422),
    .S1(net429),
    .X(_03842_));
 sky130_fd_sc_hd__mux4_2 _27141_ (.A0(_03839_),
    .A1(_03840_),
    .A2(_03841_),
    .A3(_03842_),
    .S0(net416),
    .S1(net414),
    .X(_03843_));
 sky130_fd_sc_hd__mux4_2 _27142_ (.A0(\w[33][1] ),
    .A1(\w[37][1] ),
    .A2(\w[35][1] ),
    .A3(\w[39][1] ),
    .S0(net422),
    .S1(net429),
    .X(_03844_));
 sky130_fd_sc_hd__mux4_2 _27143_ (.A0(\w[41][1] ),
    .A1(\w[45][1] ),
    .A2(\w[43][1] ),
    .A3(\w[47][1] ),
    .S0(net424),
    .S1(net429),
    .X(_03845_));
 sky130_fd_sc_hd__mux4_2 _27144_ (.A0(\w[49][1] ),
    .A1(\w[53][1] ),
    .A2(\w[51][1] ),
    .A3(\w[55][1] ),
    .S0(net422),
    .S1(net429),
    .X(_03846_));
 sky130_fd_sc_hd__mux4_2 _27145_ (.A0(\w[57][1] ),
    .A1(\w[61][1] ),
    .A2(\w[59][1] ),
    .A3(\w[63][1] ),
    .S0(net424),
    .S1(net429),
    .X(_03847_));
 sky130_fd_sc_hd__mux4_2 _27146_ (.A0(_03844_),
    .A1(_03845_),
    .A2(_03846_),
    .A3(_03847_),
    .S0(net417),
    .S1(net540),
    .X(_03848_));
 sky130_fd_sc_hd__mux2i_4 _27147_ (.A0(_03843_),
    .A1(_03848_),
    .S(net413),
    .Y(_03849_));
 sky130_fd_sc_hd__xnor2_1 _27148_ (.A(_03743_),
    .B(_03849_),
    .Y(_03850_));
 sky130_fd_sc_hd__xnor2_1 _27149_ (.A(_03320_),
    .B(_03850_),
    .Y(_11941_));
 sky130_fd_sc_hd__mux4_2 _27150_ (.A0(\w[0][0] ),
    .A1(\w[4][0] ),
    .A2(\w[2][0] ),
    .A3(\w[6][0] ),
    .S0(net500),
    .S1(net507),
    .X(_03851_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_4 ();
 sky130_fd_sc_hd__mux4_2 _27152_ (.A0(\w[8][0] ),
    .A1(\w[12][0] ),
    .A2(\w[10][0] ),
    .A3(\w[14][0] ),
    .S0(net500),
    .S1(net507),
    .X(_03853_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_2 ();
 sky130_fd_sc_hd__mux4_2 _27155_ (.A0(\w[16][0] ),
    .A1(\w[20][0] ),
    .A2(\w[18][0] ),
    .A3(\w[22][0] ),
    .S0(net500),
    .S1(net507),
    .X(_03856_));
 sky130_fd_sc_hd__mux4_2 _27156_ (.A0(\w[24][0] ),
    .A1(\w[28][0] ),
    .A2(\w[26][0] ),
    .A3(\w[30][0] ),
    .S0(net500),
    .S1(net507),
    .X(_03857_));
 sky130_fd_sc_hd__mux4_2 _27157_ (.A0(_03851_),
    .A1(_03853_),
    .A2(_03856_),
    .A3(_03857_),
    .S0(net497),
    .S1(net495),
    .X(_03858_));
 sky130_fd_sc_hd__mux4_2 _27158_ (.A0(\w[32][0] ),
    .A1(\w[36][0] ),
    .A2(\w[34][0] ),
    .A3(\w[38][0] ),
    .S0(net502),
    .S1(net508),
    .X(_03859_));
 sky130_fd_sc_hd__mux4_2 _27159_ (.A0(\w[40][0] ),
    .A1(\w[44][0] ),
    .A2(\w[42][0] ),
    .A3(\w[46][0] ),
    .S0(net502),
    .S1(net508),
    .X(_03860_));
 sky130_fd_sc_hd__mux4_2 _27160_ (.A0(\w[48][0] ),
    .A1(\w[52][0] ),
    .A2(\w[50][0] ),
    .A3(\w[54][0] ),
    .S0(net502),
    .S1(net508),
    .X(_03861_));
 sky130_fd_sc_hd__mux4_2 _27161_ (.A0(\w[56][0] ),
    .A1(\w[60][0] ),
    .A2(\w[58][0] ),
    .A3(\w[62][0] ),
    .S0(net502),
    .S1(net508),
    .X(_03862_));
 sky130_fd_sc_hd__mux4_2 _27162_ (.A0(_03859_),
    .A1(_03860_),
    .A2(_03861_),
    .A3(_03862_),
    .S0(net497),
    .S1(net495),
    .X(_03863_));
 sky130_fd_sc_hd__mux2i_4 _27163_ (.A0(_03858_),
    .A1(_03863_),
    .S(net492),
    .Y(_03864_));
 sky130_fd_sc_hd__xnor2_1 _27164_ (.A(_03656_),
    .B(_03864_),
    .Y(_03865_));
 sky130_fd_sc_hd__xnor2_1 _27165_ (.A(_03181_),
    .B(_03865_),
    .Y(_11940_));
 sky130_fd_sc_hd__mux4_2 _27166_ (.A0(\w[0][14] ),
    .A1(\w[4][14] ),
    .A2(\w[2][14] ),
    .A3(\w[6][14] ),
    .S0(net386),
    .S1(net393),
    .X(_03866_));
 sky130_fd_sc_hd__mux4_2 _27167_ (.A0(\w[8][14] ),
    .A1(\w[12][14] ),
    .A2(\w[10][14] ),
    .A3(\w[14][14] ),
    .S0(net386),
    .S1(net393),
    .X(_03867_));
 sky130_fd_sc_hd__mux4_2 _27168_ (.A0(\w[16][14] ),
    .A1(\w[20][14] ),
    .A2(\w[18][14] ),
    .A3(\w[22][14] ),
    .S0(net386),
    .S1(net393),
    .X(_03868_));
 sky130_fd_sc_hd__mux4_2 _27169_ (.A0(\w[24][14] ),
    .A1(\w[28][14] ),
    .A2(\w[26][14] ),
    .A3(\w[30][14] ),
    .S0(net386),
    .S1(net393),
    .X(_03869_));
 sky130_fd_sc_hd__mux4_2 _27170_ (.A0(_03866_),
    .A1(_03867_),
    .A2(_03868_),
    .A3(_03869_),
    .S0(net377),
    .S1(net375),
    .X(_03870_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_1 ();
 sky130_fd_sc_hd__mux4_2 _27172_ (.A0(\w[32][14] ),
    .A1(\w[36][14] ),
    .A2(\w[34][14] ),
    .A3(\w[38][14] ),
    .S0(net385),
    .S1(net392),
    .X(_03872_));
 sky130_fd_sc_hd__mux4_2 _27173_ (.A0(\w[40][14] ),
    .A1(\w[44][14] ),
    .A2(\w[42][14] ),
    .A3(\w[46][14] ),
    .S0(net385),
    .S1(net392),
    .X(_03873_));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_0 ();
 sky130_fd_sc_hd__mux4_2 _27175_ (.A0(\w[48][14] ),
    .A1(\w[52][14] ),
    .A2(\w[50][14] ),
    .A3(\w[54][14] ),
    .S0(net385),
    .S1(net392),
    .X(_03875_));
 sky130_fd_sc_hd__mux4_2 _27176_ (.A0(\w[56][14] ),
    .A1(\w[60][14] ),
    .A2(\w[58][14] ),
    .A3(\w[62][14] ),
    .S0(net385),
    .S1(net392),
    .X(_03876_));
 sky130_fd_sc_hd__mux4_2 _27177_ (.A0(_03872_),
    .A1(_03873_),
    .A2(_03875_),
    .A3(_03876_),
    .S0(net377),
    .S1(net375),
    .X(_03877_));
 sky130_fd_sc_hd__mux2i_4 _27178_ (.A0(_03870_),
    .A1(_03877_),
    .S(net373),
    .Y(_11939_));
 sky130_fd_sc_hd__mux4_2 _27179_ (.A0(\w[1][14] ),
    .A1(\w[5][14] ),
    .A2(\w[3][14] ),
    .A3(\w[7][14] ),
    .S0(net464),
    .S1(net468),
    .X(_03878_));
 sky130_fd_sc_hd__mux4_2 _27180_ (.A0(\w[9][14] ),
    .A1(\w[13][14] ),
    .A2(\w[11][14] ),
    .A3(\w[15][14] ),
    .S0(net464),
    .S1(net468),
    .X(_03879_));
 sky130_fd_sc_hd__mux4_2 _27181_ (.A0(\w[17][14] ),
    .A1(\w[21][14] ),
    .A2(\w[19][14] ),
    .A3(\w[23][14] ),
    .S0(net464),
    .S1(net468),
    .X(_03880_));
 sky130_fd_sc_hd__mux4_2 _27182_ (.A0(\w[25][14] ),
    .A1(\w[29][14] ),
    .A2(\w[27][14] ),
    .A3(\w[31][14] ),
    .S0(net464),
    .S1(net468),
    .X(_03881_));
 sky130_fd_sc_hd__mux4_2 _27183_ (.A0(_03878_),
    .A1(_03879_),
    .A2(_03880_),
    .A3(_03881_),
    .S0(\count16_2[3] ),
    .S1(net454),
    .X(_03882_));
 sky130_fd_sc_hd__fa_1 _27184_ (.A(_11579_),
    .B(_11580_),
    .CIN(_11581_),
    .COUT(_11582_),
    .SUM(_11583_));
 sky130_fd_sc_hd__fa_1 _27185_ (.A(_11584_),
    .B(_11585_),
    .CIN(_11586_),
    .COUT(_11587_),
    .SUM(_11588_));
 sky130_fd_sc_hd__fa_1 _27186_ (.A(_11589_),
    .B(_11582_),
    .CIN(_11588_),
    .COUT(_11590_),
    .SUM(_11591_));
 sky130_fd_sc_hd__fa_1 _27187_ (.A(_11592_),
    .B(_11593_),
    .CIN(_11594_),
    .COUT(_11595_),
    .SUM(_11596_));
 sky130_fd_sc_hd__fa_1 _27188_ (.A(_11597_),
    .B(_11587_),
    .CIN(_11596_),
    .COUT(_11598_),
    .SUM(_11599_));
 sky130_fd_sc_hd__fa_1 _27189_ (.A(_11600_),
    .B(_11590_),
    .CIN(_11599_),
    .COUT(_11601_),
    .SUM(_11602_));
 sky130_fd_sc_hd__fa_1 _27190_ (.A(_11603_),
    .B(_11604_),
    .CIN(_11605_),
    .COUT(_11606_),
    .SUM(_11607_));
 sky130_fd_sc_hd__fa_1 _27191_ (.A(_11608_),
    .B(_11595_),
    .CIN(_11607_),
    .COUT(_11609_),
    .SUM(_11610_));
 sky130_fd_sc_hd__fa_1 _27192_ (.A(_11611_),
    .B(_11612_),
    .CIN(_11613_),
    .COUT(_11614_),
    .SUM(_11615_));
 sky130_fd_sc_hd__fa_1 _27193_ (.A(_11616_),
    .B(_11606_),
    .CIN(_11615_),
    .COUT(_11617_),
    .SUM(_11618_));
 sky130_fd_sc_hd__fa_1 _27194_ (.A(_11619_),
    .B(_11620_),
    .CIN(_11621_),
    .COUT(_11622_),
    .SUM(_11623_));
 sky130_fd_sc_hd__fa_1 _27195_ (.A(_11624_),
    .B(_11614_),
    .CIN(_11623_),
    .COUT(_11625_),
    .SUM(_11626_));
 sky130_fd_sc_hd__fa_1 _27196_ (.A(_11627_),
    .B(_11628_),
    .CIN(_11629_),
    .COUT(_11630_),
    .SUM(_11631_));
 sky130_fd_sc_hd__fa_1 _27197_ (.A(_11632_),
    .B(_11622_),
    .CIN(_11631_),
    .COUT(_11633_),
    .SUM(_11634_));
 sky130_fd_sc_hd__fa_1 _27198_ (.A(_11635_),
    .B(_11636_),
    .CIN(_11637_),
    .COUT(_11638_),
    .SUM(_11639_));
 sky130_fd_sc_hd__fa_1 _27199_ (.A(_11640_),
    .B(_11630_),
    .CIN(_11639_),
    .COUT(_11641_),
    .SUM(_11642_));
 sky130_fd_sc_hd__fa_1 _27200_ (.A(_11643_),
    .B(_11644_),
    .CIN(_11645_),
    .COUT(_11646_),
    .SUM(_11647_));
 sky130_fd_sc_hd__fa_1 _27201_ (.A(_11648_),
    .B(_11638_),
    .CIN(_11647_),
    .COUT(_11649_),
    .SUM(_11650_));
 sky130_fd_sc_hd__fa_1 _27202_ (.A(_11651_),
    .B(_11652_),
    .CIN(_11653_),
    .COUT(_11654_),
    .SUM(_11655_));
 sky130_fd_sc_hd__fa_1 _27203_ (.A(_11656_),
    .B(_11646_),
    .CIN(_11655_),
    .COUT(_11657_),
    .SUM(_11658_));
 sky130_fd_sc_hd__fa_1 _27204_ (.A(_11659_),
    .B(_11660_),
    .CIN(_11661_),
    .COUT(_11662_),
    .SUM(_11663_));
 sky130_fd_sc_hd__fa_1 _27205_ (.A(_11664_),
    .B(_11654_),
    .CIN(_11663_),
    .COUT(_11665_),
    .SUM(_11666_));
 sky130_fd_sc_hd__fa_1 _27206_ (.A(_11667_),
    .B(_11668_),
    .CIN(_11669_),
    .COUT(_11670_),
    .SUM(_11671_));
 sky130_fd_sc_hd__fa_1 _27207_ (.A(_11672_),
    .B(_11662_),
    .CIN(_11671_),
    .COUT(_11673_),
    .SUM(_11674_));
 sky130_fd_sc_hd__fa_1 _27208_ (.A(_11675_),
    .B(_11676_),
    .CIN(_11677_),
    .COUT(_11678_),
    .SUM(_11679_));
 sky130_fd_sc_hd__fa_1 _27209_ (.A(_11680_),
    .B(_11670_),
    .CIN(_11679_),
    .COUT(_11681_),
    .SUM(_11682_));
 sky130_fd_sc_hd__fa_1 _27210_ (.A(_11683_),
    .B(_11684_),
    .CIN(_11685_),
    .COUT(_11686_),
    .SUM(_11687_));
 sky130_fd_sc_hd__fa_1 _27211_ (.A(_11688_),
    .B(_11678_),
    .CIN(_11687_),
    .COUT(_11689_),
    .SUM(_11690_));
 sky130_fd_sc_hd__fa_1 _27212_ (.A(_11691_),
    .B(_11692_),
    .CIN(_11693_),
    .COUT(_11694_),
    .SUM(_11695_));
 sky130_fd_sc_hd__fa_1 _27213_ (.A(_11696_),
    .B(_11686_),
    .CIN(_11695_),
    .COUT(_11697_),
    .SUM(_11698_));
 sky130_fd_sc_hd__fa_1 _27214_ (.A(_11699_),
    .B(_11700_),
    .CIN(_11701_),
    .COUT(_11702_),
    .SUM(_11703_));
 sky130_fd_sc_hd__fa_1 _27215_ (.A(_11704_),
    .B(_11694_),
    .CIN(_11703_),
    .COUT(_11705_),
    .SUM(_11706_));
 sky130_fd_sc_hd__fa_1 _27216_ (.A(_11707_),
    .B(_11708_),
    .CIN(_11709_),
    .COUT(_11710_),
    .SUM(_11711_));
 sky130_fd_sc_hd__fa_1 _27217_ (.A(_11712_),
    .B(_11702_),
    .CIN(_11711_),
    .COUT(_11713_),
    .SUM(_11714_));
 sky130_fd_sc_hd__fa_1 _27218_ (.A(_11715_),
    .B(_11716_),
    .CIN(_11717_),
    .COUT(_11718_),
    .SUM(_11719_));
 sky130_fd_sc_hd__fa_1 _27219_ (.A(_11720_),
    .B(_11710_),
    .CIN(_11719_),
    .COUT(_11721_),
    .SUM(_11722_));
 sky130_fd_sc_hd__fa_1 _27220_ (.A(_11723_),
    .B(_11724_),
    .CIN(_11725_),
    .COUT(_11726_),
    .SUM(_11727_));
 sky130_fd_sc_hd__fa_1 _27221_ (.A(_11728_),
    .B(_11718_),
    .CIN(_11727_),
    .COUT(_11729_),
    .SUM(_11730_));
 sky130_fd_sc_hd__fa_1 _27222_ (.A(_11731_),
    .B(_11732_),
    .CIN(_11733_),
    .COUT(_11734_),
    .SUM(_11735_));
 sky130_fd_sc_hd__fa_1 _27223_ (.A(_11736_),
    .B(_11726_),
    .CIN(_11735_),
    .COUT(_11737_),
    .SUM(_11738_));
 sky130_fd_sc_hd__fa_1 _27224_ (.A(_11739_),
    .B(_11740_),
    .CIN(_11741_),
    .COUT(_11742_),
    .SUM(_11743_));
 sky130_fd_sc_hd__fa_1 _27225_ (.A(_11744_),
    .B(_11734_),
    .CIN(_11743_),
    .COUT(_11745_),
    .SUM(_11746_));
 sky130_fd_sc_hd__fa_1 _27226_ (.A(_11747_),
    .B(_11748_),
    .CIN(_11749_),
    .COUT(_11750_),
    .SUM(_11751_));
 sky130_fd_sc_hd__fa_1 _27227_ (.A(_11752_),
    .B(_11742_),
    .CIN(_11751_),
    .COUT(_11753_),
    .SUM(_11754_));
 sky130_fd_sc_hd__fa_1 _27228_ (.A(_11755_),
    .B(_11756_),
    .CIN(_11757_),
    .COUT(_11758_),
    .SUM(_11759_));
 sky130_fd_sc_hd__fa_1 _27229_ (.A(_11760_),
    .B(_11750_),
    .CIN(_11759_),
    .COUT(_11761_),
    .SUM(_11762_));
 sky130_fd_sc_hd__fa_1 _27230_ (.A(_11763_),
    .B(_11764_),
    .CIN(_11765_),
    .COUT(_11766_),
    .SUM(_11767_));
 sky130_fd_sc_hd__fa_1 _27231_ (.A(_11768_),
    .B(_11758_),
    .CIN(_11767_),
    .COUT(_11769_),
    .SUM(_11770_));
 sky130_fd_sc_hd__fa_1 _27232_ (.A(_11771_),
    .B(_11772_),
    .CIN(_11773_),
    .COUT(_11774_),
    .SUM(_11775_));
 sky130_fd_sc_hd__fa_1 _27233_ (.A(_11776_),
    .B(_11766_),
    .CIN(_11775_),
    .COUT(_11777_),
    .SUM(_11778_));
 sky130_fd_sc_hd__fa_1 _27234_ (.A(_11779_),
    .B(_11780_),
    .CIN(_11781_),
    .COUT(_11782_),
    .SUM(_11783_));
 sky130_fd_sc_hd__fa_1 _27235_ (.A(_11784_),
    .B(_11774_),
    .CIN(_11783_),
    .COUT(_11785_),
    .SUM(_11786_));
 sky130_fd_sc_hd__fa_1 _27236_ (.A(_11787_),
    .B(_11788_),
    .CIN(_11789_),
    .COUT(_11790_),
    .SUM(_11791_));
 sky130_fd_sc_hd__fa_1 _27237_ (.A(_11792_),
    .B(_11782_),
    .CIN(_11791_),
    .COUT(_11793_),
    .SUM(_11794_));
 sky130_fd_sc_hd__fa_1 _27238_ (.A(_11795_),
    .B(_11796_),
    .CIN(_11797_),
    .COUT(_11798_),
    .SUM(_11799_));
 sky130_fd_sc_hd__fa_1 _27239_ (.A(_11800_),
    .B(_11790_),
    .CIN(_11799_),
    .COUT(_11801_),
    .SUM(_11802_));
 sky130_fd_sc_hd__fa_1 _27240_ (.A(_11803_),
    .B(_11804_),
    .CIN(_11805_),
    .COUT(_11806_),
    .SUM(_11807_));
 sky130_fd_sc_hd__fa_1 _27241_ (.A(_11808_),
    .B(_11798_),
    .CIN(_11807_),
    .COUT(_11809_),
    .SUM(_11810_));
 sky130_fd_sc_hd__fa_1 _27242_ (.A(_11811_),
    .B(_11812_),
    .CIN(_11813_),
    .COUT(_11814_),
    .SUM(_11815_));
 sky130_fd_sc_hd__fa_1 _27243_ (.A(_11816_),
    .B(_11806_),
    .CIN(_11815_),
    .COUT(_11817_),
    .SUM(_11818_));
 sky130_fd_sc_hd__fa_1 _27244_ (.A(_11819_),
    .B(_11820_),
    .CIN(_11821_),
    .COUT(_11822_),
    .SUM(_11823_));
 sky130_fd_sc_hd__fa_1 _27245_ (.A(_11824_),
    .B(_11814_),
    .CIN(_11823_),
    .COUT(_11825_),
    .SUM(_11826_));
 sky130_fd_sc_hd__fa_1 _27246_ (.A(_11827_),
    .B(_11828_),
    .CIN(_11829_),
    .COUT(_11830_),
    .SUM(_11831_));
 sky130_fd_sc_hd__fa_1 _27247_ (.A(_11832_),
    .B(_11833_),
    .CIN(_11834_),
    .COUT(_11835_),
    .SUM(_11836_));
 sky130_fd_sc_hd__fa_1 _27248_ (.A(_11837_),
    .B(_11830_),
    .CIN(_11836_),
    .COUT(_11838_),
    .SUM(_11839_));
 sky130_fd_sc_hd__fa_1 _27249_ (.A(_11840_),
    .B(_11841_),
    .CIN(_11842_),
    .COUT(_11843_),
    .SUM(_11844_));
 sky130_fd_sc_hd__fa_1 _27250_ (.A(_11845_),
    .B(_11835_),
    .CIN(_11844_),
    .COUT(_11846_),
    .SUM(_11847_));
 sky130_fd_sc_hd__fa_1 _27251_ (.A(_11848_),
    .B(_11838_),
    .CIN(_11847_),
    .COUT(_11849_),
    .SUM(_11850_));
 sky130_fd_sc_hd__fa_1 _27252_ (.A(_11851_),
    .B(_11852_),
    .CIN(_11853_),
    .COUT(_11854_),
    .SUM(_11855_));
 sky130_fd_sc_hd__fa_1 _27253_ (.A(_11856_),
    .B(_11843_),
    .CIN(_11855_),
    .COUT(_11857_),
    .SUM(_11858_));
 sky130_fd_sc_hd__fa_1 _27254_ (.A(_11859_),
    .B(_11860_),
    .CIN(_11861_),
    .COUT(_11862_),
    .SUM(_11863_));
 sky130_fd_sc_hd__fa_1 _27255_ (.A(_11864_),
    .B(_11854_),
    .CIN(_11863_),
    .COUT(_11865_),
    .SUM(_11866_));
 sky130_fd_sc_hd__fa_1 _27256_ (.A(_11867_),
    .B(_11868_),
    .CIN(_11869_),
    .COUT(_11870_),
    .SUM(_11871_));
 sky130_fd_sc_hd__fa_1 _27257_ (.A(_11872_),
    .B(_11862_),
    .CIN(_11871_),
    .COUT(_11873_),
    .SUM(_11874_));
 sky130_fd_sc_hd__fa_1 _27258_ (.A(_11875_),
    .B(_11876_),
    .CIN(_11877_),
    .COUT(_11878_),
    .SUM(_11879_));
 sky130_fd_sc_hd__fa_1 _27259_ (.A(_11880_),
    .B(_11870_),
    .CIN(_11879_),
    .COUT(_11881_),
    .SUM(_11882_));
 sky130_fd_sc_hd__fa_1 _27260_ (.A(_11883_),
    .B(_11884_),
    .CIN(_11885_),
    .COUT(_11886_),
    .SUM(_11887_));
 sky130_fd_sc_hd__fa_1 _27261_ (.A(_11888_),
    .B(_11878_),
    .CIN(_11887_),
    .COUT(_11889_),
    .SUM(_11890_));
 sky130_fd_sc_hd__fa_1 _27262_ (.A(_11891_),
    .B(_11892_),
    .CIN(_11893_),
    .COUT(_11894_),
    .SUM(_11895_));
 sky130_fd_sc_hd__fa_1 _27263_ (.A(_11896_),
    .B(_11886_),
    .CIN(_11895_),
    .COUT(_11897_),
    .SUM(_11898_));
 sky130_fd_sc_hd__fa_1 _27264_ (.A(_11899_),
    .B(_11900_),
    .CIN(_11901_),
    .COUT(_11902_),
    .SUM(_11903_));
 sky130_fd_sc_hd__fa_1 _27265_ (.A(_11904_),
    .B(_11894_),
    .CIN(_11903_),
    .COUT(_11905_),
    .SUM(_11906_));
 sky130_fd_sc_hd__fa_1 _27266_ (.A(_11907_),
    .B(_11908_),
    .CIN(_11909_),
    .COUT(_11910_),
    .SUM(_11911_));
 sky130_fd_sc_hd__fa_1 _27267_ (.A(_11912_),
    .B(_11902_),
    .CIN(_11911_),
    .COUT(_11913_),
    .SUM(_11914_));
 sky130_fd_sc_hd__fa_1 _27268_ (.A(_11915_),
    .B(_11916_),
    .CIN(_11917_),
    .COUT(_11918_),
    .SUM(_11919_));
 sky130_fd_sc_hd__fa_1 _27269_ (.A(_11920_),
    .B(_11910_),
    .CIN(_11919_),
    .COUT(_11921_),
    .SUM(_11922_));
 sky130_fd_sc_hd__fa_1 _27270_ (.A(_11923_),
    .B(_11924_),
    .CIN(_11925_),
    .COUT(_11926_),
    .SUM(_11927_));
 sky130_fd_sc_hd__fa_1 _27271_ (.A(_11928_),
    .B(_11918_),
    .CIN(_11927_),
    .COUT(_11929_),
    .SUM(_11930_));
 sky130_fd_sc_hd__fa_1 _27272_ (.A(_11931_),
    .B(_11932_),
    .CIN(_11933_),
    .COUT(_11934_),
    .SUM(_11935_));
 sky130_fd_sc_hd__fa_1 _27273_ (.A(_11936_),
    .B(_11926_),
    .CIN(_11935_),
    .COUT(_11937_),
    .SUM(_11938_));
 sky130_fd_sc_hd__fa_1 _27274_ (.A(_11939_),
    .B(_11940_),
    .CIN(_11941_),
    .COUT(_11942_),
    .SUM(_11943_));
 sky130_fd_sc_hd__fa_1 _27275_ (.A(_11944_),
    .B(_11934_),
    .CIN(_11943_),
    .COUT(_11945_),
    .SUM(_11946_));
 sky130_fd_sc_hd__fa_1 _27276_ (.A(_11947_),
    .B(_11948_),
    .CIN(_11949_),
    .COUT(_11950_),
    .SUM(_11951_));
 sky130_fd_sc_hd__fa_1 _27277_ (.A(_11952_),
    .B(_11942_),
    .CIN(_11951_),
    .COUT(_11953_),
    .SUM(_11954_));
 sky130_fd_sc_hd__fa_1 _27278_ (.A(_11955_),
    .B(_11956_),
    .CIN(_11957_),
    .COUT(_11958_),
    .SUM(_11959_));
 sky130_fd_sc_hd__fa_1 _27279_ (.A(_11960_),
    .B(_11950_),
    .CIN(_11959_),
    .COUT(_11961_),
    .SUM(_11962_));
 sky130_fd_sc_hd__fa_1 _27280_ (.A(_11963_),
    .B(_11964_),
    .CIN(_11965_),
    .COUT(_11966_),
    .SUM(_11967_));
 sky130_fd_sc_hd__fa_1 _27281_ (.A(_11968_),
    .B(_11958_),
    .CIN(_11967_),
    .COUT(_11969_),
    .SUM(_11970_));
 sky130_fd_sc_hd__fa_1 _27282_ (.A(_11971_),
    .B(_11972_),
    .CIN(_11973_),
    .COUT(_11974_),
    .SUM(_11975_));
 sky130_fd_sc_hd__fa_1 _27283_ (.A(_11976_),
    .B(_11966_),
    .CIN(_11975_),
    .COUT(_11977_),
    .SUM(_11978_));
 sky130_fd_sc_hd__fa_1 _27284_ (.A(_11979_),
    .B(_11980_),
    .CIN(_11981_),
    .COUT(_11982_),
    .SUM(_11983_));
 sky130_fd_sc_hd__fa_1 _27285_ (.A(_11984_),
    .B(_11974_),
    .CIN(_11983_),
    .COUT(_11985_),
    .SUM(_11986_));
 sky130_fd_sc_hd__fa_1 _27286_ (.A(_11987_),
    .B(_11988_),
    .CIN(_11989_),
    .COUT(_11990_),
    .SUM(_11991_));
 sky130_fd_sc_hd__fa_1 _27287_ (.A(_11992_),
    .B(_11982_),
    .CIN(_11991_),
    .COUT(_11993_),
    .SUM(_11994_));
 sky130_fd_sc_hd__fa_1 _27288_ (.A(_11995_),
    .B(_11996_),
    .CIN(_11997_),
    .COUT(_11998_),
    .SUM(_11999_));
 sky130_fd_sc_hd__fa_1 _27289_ (.A(_12000_),
    .B(_11990_),
    .CIN(_11999_),
    .COUT(_12001_),
    .SUM(_12002_));
 sky130_fd_sc_hd__fa_1 _27290_ (.A(_12003_),
    .B(_12004_),
    .CIN(_12005_),
    .COUT(_12006_),
    .SUM(_12007_));
 sky130_fd_sc_hd__fa_1 _27291_ (.A(_12008_),
    .B(_11998_),
    .CIN(_12007_),
    .COUT(_12009_),
    .SUM(_12010_));
 sky130_fd_sc_hd__fa_1 _27292_ (.A(_12011_),
    .B(_12012_),
    .CIN(_12013_),
    .COUT(_12014_),
    .SUM(_12015_));
 sky130_fd_sc_hd__fa_1 _27293_ (.A(_12016_),
    .B(_12006_),
    .CIN(_12015_),
    .COUT(_12017_),
    .SUM(_12018_));
 sky130_fd_sc_hd__fa_1 _27294_ (.A(_12019_),
    .B(_12020_),
    .CIN(_12021_),
    .COUT(_12022_),
    .SUM(_12023_));
 sky130_fd_sc_hd__fa_1 _27295_ (.A(_12024_),
    .B(_12014_),
    .CIN(_12023_),
    .COUT(_12025_),
    .SUM(_12026_));
 sky130_fd_sc_hd__fa_1 _27296_ (.A(_12027_),
    .B(_12028_),
    .CIN(_12029_),
    .COUT(_12030_),
    .SUM(_12031_));
 sky130_fd_sc_hd__fa_1 _27297_ (.A(_12032_),
    .B(_12022_),
    .CIN(_12031_),
    .COUT(_12033_),
    .SUM(_12034_));
 sky130_fd_sc_hd__fa_1 _27298_ (.A(_12035_),
    .B(_12036_),
    .CIN(_12037_),
    .COUT(_12038_),
    .SUM(_12039_));
 sky130_fd_sc_hd__fa_1 _27299_ (.A(_12040_),
    .B(_12030_),
    .CIN(_12039_),
    .COUT(_12041_),
    .SUM(_12042_));
 sky130_fd_sc_hd__fa_1 _27300_ (.A(_12043_),
    .B(_12044_),
    .CIN(_12045_),
    .COUT(_12046_),
    .SUM(_12047_));
 sky130_fd_sc_hd__fa_1 _27301_ (.A(_12048_),
    .B(_12038_),
    .CIN(_12047_),
    .COUT(_12049_),
    .SUM(_12050_));
 sky130_fd_sc_hd__fa_1 _27302_ (.A(_12051_),
    .B(_12052_),
    .CIN(_12053_),
    .COUT(_12054_),
    .SUM(_12055_));
 sky130_fd_sc_hd__fa_1 _27303_ (.A(_12056_),
    .B(_12046_),
    .CIN(_12055_),
    .COUT(_12057_),
    .SUM(_12058_));
 sky130_fd_sc_hd__fa_1 _27304_ (.A(_12059_),
    .B(_12060_),
    .CIN(_12061_),
    .COUT(_12062_),
    .SUM(_12063_));
 sky130_fd_sc_hd__fa_1 _27305_ (.A(_12064_),
    .B(_12054_),
    .CIN(_12063_),
    .COUT(_12065_),
    .SUM(_12066_));
 sky130_fd_sc_hd__fa_1 _27306_ (.A(_12067_),
    .B(_12068_),
    .CIN(_12069_),
    .COUT(_12070_),
    .SUM(_12071_));
 sky130_fd_sc_hd__fa_1 _27307_ (.A(_12072_),
    .B(_12062_),
    .CIN(_12071_),
    .COUT(_12073_),
    .SUM(_12074_));
 sky130_fd_sc_hd__fa_1 _27308_ (.A(_12075_),
    .B(_12076_),
    .CIN(_12077_),
    .COUT(_12078_),
    .SUM(_12079_));
 sky130_fd_sc_hd__fa_2 _27309_ (.A(\hash.CA2.p1[1] ),
    .B(\hash.CA2.p3[1] ),
    .CIN(_12080_),
    .COUT(_12081_),
    .SUM(_12082_));
 sky130_fd_sc_hd__fa_2 _27310_ (.A(_12085_),
    .B(_12084_),
    .CIN(_12083_),
    .COUT(_12086_),
    .SUM(_12087_));
 sky130_fd_sc_hd__fa_1 _27311_ (.A(_12087_),
    .B(_12088_),
    .CIN(_12089_),
    .COUT(_12090_),
    .SUM(_12091_));
 sky130_fd_sc_hd__fa_1 _27312_ (.A(\hash.CA2.p4[1] ),
    .B(_12092_),
    .CIN(_12093_),
    .COUT(_12094_),
    .SUM(_12095_));
 sky130_fd_sc_hd__fa_1 _27313_ (.A(_12096_),
    .B(_12097_),
    .CIN(_12098_),
    .COUT(_12099_),
    .SUM(_12100_));
 sky130_fd_sc_hd__fa_1 _27314_ (.A(\hash.CA2.p4[2] ),
    .B(_12101_),
    .CIN(_12102_),
    .COUT(_12103_),
    .SUM(_12104_));
 sky130_fd_sc_hd__fa_2 _27315_ (.A(_12105_),
    .B(_12106_),
    .CIN(_12107_),
    .COUT(_12108_),
    .SUM(_12109_));
 sky130_fd_sc_hd__fa_1 _27316_ (.A(_12110_),
    .B(_12111_),
    .CIN(_12112_),
    .COUT(_12113_),
    .SUM(_12114_));
 sky130_fd_sc_hd__fa_1 _27317_ (.A(\hash.CA2.p4[3] ),
    .B(_12115_),
    .CIN(_12116_),
    .COUT(_12117_),
    .SUM(_12118_));
 sky130_fd_sc_hd__fa_1 _27318_ (.A(_12119_),
    .B(_12120_),
    .CIN(_12121_),
    .COUT(_12122_),
    .SUM(_12123_));
 sky130_fd_sc_hd__fa_1 _27319_ (.A(\hash.CA2.p4[4] ),
    .B(_12124_),
    .CIN(_12125_),
    .COUT(_12126_),
    .SUM(_12127_));
 sky130_fd_sc_hd__fa_1 _27320_ (.A(_12128_),
    .B(_12129_),
    .CIN(_12130_),
    .COUT(_12131_),
    .SUM(_12132_));
 sky130_fd_sc_hd__fa_1 _27321_ (.A(\hash.CA2.p4[5] ),
    .B(_12133_),
    .CIN(_12134_),
    .COUT(_12135_),
    .SUM(_12136_));
 sky130_fd_sc_hd__fa_1 _27322_ (.A(_12137_),
    .B(_12138_),
    .CIN(_12139_),
    .COUT(_12140_),
    .SUM(_12141_));
 sky130_fd_sc_hd__fa_1 _27323_ (.A(\hash.CA2.p4[6] ),
    .B(_12142_),
    .CIN(_12143_),
    .COUT(_12144_),
    .SUM(_12145_));
 sky130_fd_sc_hd__fa_1 _27324_ (.A(_12146_),
    .B(_12147_),
    .CIN(_12148_),
    .COUT(_12149_),
    .SUM(_12150_));
 sky130_fd_sc_hd__fa_1 _27325_ (.A(\hash.CA2.p4[7] ),
    .B(_12151_),
    .CIN(_12152_),
    .COUT(_12153_),
    .SUM(_12154_));
 sky130_fd_sc_hd__fa_1 _27326_ (.A(_12157_),
    .B(_12156_),
    .CIN(_12155_),
    .COUT(_12158_),
    .SUM(_12159_));
 sky130_fd_sc_hd__fa_1 _27327_ (.A(\hash.CA2.p4[8] ),
    .B(_12160_),
    .CIN(_12161_),
    .COUT(_12162_),
    .SUM(_12163_));
 sky130_fd_sc_hd__fa_1 _27328_ (.A(_12164_),
    .B(_12165_),
    .CIN(_12166_),
    .COUT(_12167_),
    .SUM(_12168_));
 sky130_fd_sc_hd__fa_1 _27329_ (.A(\hash.CA2.p4[9] ),
    .B(_12169_),
    .CIN(_12170_),
    .COUT(_12171_),
    .SUM(_12172_));
 sky130_fd_sc_hd__fa_1 _27330_ (.A(_12173_),
    .B(_12174_),
    .CIN(_12175_),
    .COUT(_12176_),
    .SUM(_12177_));
 sky130_fd_sc_hd__fa_1 _27331_ (.A(\hash.CA2.p4[10] ),
    .B(_12178_),
    .CIN(_12179_),
    .COUT(_12180_),
    .SUM(_12181_));
 sky130_fd_sc_hd__fa_1 _27332_ (.A(_12182_),
    .B(_12183_),
    .CIN(_12184_),
    .COUT(_12185_),
    .SUM(_12186_));
 sky130_fd_sc_hd__fa_1 _27333_ (.A(\hash.CA2.p4[11] ),
    .B(_12187_),
    .CIN(_12188_),
    .COUT(_12189_),
    .SUM(_12190_));
 sky130_fd_sc_hd__fa_1 _27334_ (.A(_12191_),
    .B(_12192_),
    .CIN(_12193_),
    .COUT(_12194_),
    .SUM(_12195_));
 sky130_fd_sc_hd__fa_1 _27335_ (.A(\hash.CA2.p4[12] ),
    .B(_12196_),
    .CIN(_12197_),
    .COUT(_12198_),
    .SUM(_12199_));
 sky130_fd_sc_hd__fa_1 _27336_ (.A(_12200_),
    .B(_12201_),
    .CIN(_12202_),
    .COUT(_12203_),
    .SUM(_12204_));
 sky130_fd_sc_hd__fa_1 _27337_ (.A(\hash.CA2.p4[13] ),
    .B(_12205_),
    .CIN(_12206_),
    .COUT(_12207_),
    .SUM(_12208_));
 sky130_fd_sc_hd__fa_1 _27338_ (.A(_12209_),
    .B(_12210_),
    .CIN(_12211_),
    .COUT(_12212_),
    .SUM(_12213_));
 sky130_fd_sc_hd__fa_1 _27339_ (.A(\hash.CA2.p4[14] ),
    .B(_12214_),
    .CIN(_12215_),
    .COUT(_12216_),
    .SUM(_12217_));
 sky130_fd_sc_hd__fa_1 _27340_ (.A(_12218_),
    .B(_12219_),
    .CIN(_12220_),
    .COUT(_12221_),
    .SUM(_12222_));
 sky130_fd_sc_hd__fa_1 _27341_ (.A(\hash.CA2.p4[15] ),
    .B(_12223_),
    .CIN(_12224_),
    .COUT(_12225_),
    .SUM(_12226_));
 sky130_fd_sc_hd__fa_1 _27342_ (.A(_12227_),
    .B(_12228_),
    .CIN(_12229_),
    .COUT(_12230_),
    .SUM(_12231_));
 sky130_fd_sc_hd__fa_1 _27343_ (.A(\hash.CA2.p4[16] ),
    .B(_12232_),
    .CIN(_12233_),
    .COUT(_12234_),
    .SUM(_12235_));
 sky130_fd_sc_hd__fa_1 _27344_ (.A(_12236_),
    .B(_12237_),
    .CIN(_12238_),
    .COUT(_12239_),
    .SUM(_12240_));
 sky130_fd_sc_hd__fa_1 _27345_ (.A(\hash.CA2.p4[17] ),
    .B(_12242_),
    .CIN(_12241_),
    .COUT(_12243_),
    .SUM(_12244_));
 sky130_fd_sc_hd__fa_1 _27346_ (.A(_12245_),
    .B(_12246_),
    .CIN(_12247_),
    .COUT(_12248_),
    .SUM(_12249_));
 sky130_fd_sc_hd__fa_1 _27347_ (.A(\hash.CA2.p4[18] ),
    .B(_12250_),
    .CIN(_12251_),
    .COUT(_12252_),
    .SUM(_12253_));
 sky130_fd_sc_hd__fa_1 _27348_ (.A(_12254_),
    .B(_12255_),
    .CIN(_12256_),
    .COUT(_12257_),
    .SUM(_12258_));
 sky130_fd_sc_hd__fa_1 _27349_ (.A(\hash.CA2.p4[19] ),
    .B(_12259_),
    .CIN(_12260_),
    .COUT(_12261_),
    .SUM(_12262_));
 sky130_fd_sc_hd__fa_1 _27350_ (.A(_12263_),
    .B(_12264_),
    .CIN(_12265_),
    .COUT(_12266_),
    .SUM(_12267_));
 sky130_fd_sc_hd__fa_1 _27351_ (.A(\hash.CA2.p4[20] ),
    .B(_12268_),
    .CIN(_12269_),
    .COUT(_12270_),
    .SUM(_12271_));
 sky130_fd_sc_hd__fa_1 _27352_ (.A(_12272_),
    .B(_12273_),
    .CIN(_12274_),
    .COUT(_12275_),
    .SUM(_12276_));
 sky130_fd_sc_hd__fa_1 _27353_ (.A(\hash.CA2.p4[21] ),
    .B(_12277_),
    .CIN(_12278_),
    .COUT(_12279_),
    .SUM(_12280_));
 sky130_fd_sc_hd__fa_1 _27354_ (.A(_12281_),
    .B(_12282_),
    .CIN(_12283_),
    .COUT(_12284_),
    .SUM(_12285_));
 sky130_fd_sc_hd__fa_1 _27355_ (.A(\hash.CA2.p4[22] ),
    .B(_12286_),
    .CIN(_12287_),
    .COUT(_12288_),
    .SUM(_12289_));
 sky130_fd_sc_hd__fa_1 _27356_ (.A(_12290_),
    .B(_12291_),
    .CIN(_12292_),
    .COUT(_12293_),
    .SUM(_12294_));
 sky130_fd_sc_hd__fa_1 _27357_ (.A(\hash.CA2.p4[23] ),
    .B(_12295_),
    .CIN(_12296_),
    .COUT(_12297_),
    .SUM(_12298_));
 sky130_fd_sc_hd__fa_1 _27358_ (.A(_12299_),
    .B(_12300_),
    .CIN(_12301_),
    .COUT(_12302_),
    .SUM(_12303_));
 sky130_fd_sc_hd__fa_1 _27359_ (.A(\hash.CA2.p4[24] ),
    .B(_12304_),
    .CIN(_12305_),
    .COUT(_12306_),
    .SUM(_12307_));
 sky130_fd_sc_hd__fa_1 _27360_ (.A(_12308_),
    .B(_12309_),
    .CIN(_12310_),
    .COUT(_12311_),
    .SUM(_12312_));
 sky130_fd_sc_hd__fa_1 _27361_ (.A(\hash.CA2.p4[25] ),
    .B(_12313_),
    .CIN(_12314_),
    .COUT(_12315_),
    .SUM(_12316_));
 sky130_fd_sc_hd__fa_1 _27362_ (.A(_12317_),
    .B(_12318_),
    .CIN(_12319_),
    .COUT(_12320_),
    .SUM(_12321_));
 sky130_fd_sc_hd__fa_1 _27363_ (.A(\hash.CA2.p4[26] ),
    .B(_12322_),
    .CIN(_12323_),
    .COUT(_12324_),
    .SUM(_12325_));
 sky130_fd_sc_hd__fa_1 _27364_ (.A(_12326_),
    .B(_12327_),
    .CIN(_12328_),
    .COUT(_12329_),
    .SUM(_12330_));
 sky130_fd_sc_hd__fa_1 _27365_ (.A(\hash.CA2.p4[27] ),
    .B(_12331_),
    .CIN(_12332_),
    .COUT(_12333_),
    .SUM(_12334_));
 sky130_fd_sc_hd__fa_1 _27366_ (.A(_12335_),
    .B(_12336_),
    .CIN(_12337_),
    .COUT(_12338_),
    .SUM(_12339_));
 sky130_fd_sc_hd__fa_1 _27367_ (.A(\hash.CA2.p4[28] ),
    .B(_12340_),
    .CIN(_12341_),
    .COUT(_12342_),
    .SUM(_12343_));
 sky130_fd_sc_hd__fa_1 _27368_ (.A(_12344_),
    .B(_12345_),
    .CIN(_12346_),
    .COUT(_12347_),
    .SUM(_12348_));
 sky130_fd_sc_hd__fa_1 _27369_ (.A(\hash.CA2.p4[29] ),
    .B(_12349_),
    .CIN(_12350_),
    .COUT(_12351_),
    .SUM(_12352_));
 sky130_fd_sc_hd__fa_1 _27370_ (.A(_12353_),
    .B(_12354_),
    .CIN(_12355_),
    .COUT(_12356_),
    .SUM(_12357_));
 sky130_fd_sc_hd__fa_1 _27371_ (.A(\hash.CA2.p4[30] ),
    .B(_12358_),
    .CIN(_12359_),
    .COUT(_12360_),
    .SUM(_12361_));
 sky130_fd_sc_hd__fa_1 _27372_ (.A(\hash.CA2.p5[1] ),
    .B(_12362_),
    .CIN(_12363_),
    .COUT(_12364_),
    .SUM(_12365_));
 sky130_fd_sc_hd__fa_1 _27373_ (.A(_12366_),
    .B(_12367_),
    .CIN(_12368_),
    .COUT(_12369_),
    .SUM(_12370_));
 sky130_fd_sc_hd__fa_1 _27374_ (.A(_12371_),
    .B(_12372_),
    .CIN(_00843_),
    .COUT(_12373_),
    .SUM(_12374_));
 sky130_fd_sc_hd__fa_1 _27375_ (.A(\hash.CA1.k_i2[2] ),
    .B(\hash.CA1.w_i2[2] ),
    .CIN(_12375_),
    .COUT(_12376_),
    .SUM(_12377_));
 sky130_fd_sc_hd__fa_1 _27376_ (.A(_12378_),
    .B(_12379_),
    .CIN(_12377_),
    .COUT(_12380_),
    .SUM(\hash.CA1.p4[2] ));
 sky130_fd_sc_hd__fa_1 _27377_ (.A(_12381_),
    .B(_12382_),
    .CIN(_12383_),
    .COUT(_12384_),
    .SUM(_12385_));
 sky130_fd_sc_hd__fa_1 _27378_ (.A(\hash.CA1.k_i2[4] ),
    .B(\hash.CA1.w_i2[4] ),
    .CIN(_12386_),
    .COUT(_12387_),
    .SUM(_12388_));
 sky130_fd_sc_hd__fa_1 _27379_ (.A(_12389_),
    .B(_12390_),
    .CIN(_12391_),
    .COUT(_12392_),
    .SUM(_12393_));
 sky130_fd_sc_hd__fa_1 _27380_ (.A(\hash.CA1.k_i2[6] ),
    .B(\hash.CA1.w_i2[6] ),
    .CIN(_12394_),
    .COUT(_12395_),
    .SUM(_12396_));
 sky130_fd_sc_hd__fa_1 _27381_ (.A(_12397_),
    .B(_12398_),
    .CIN(_12399_),
    .COUT(_12400_),
    .SUM(_12401_));
 sky130_fd_sc_hd__fa_1 _27382_ (.A(_12402_),
    .B(_12403_),
    .CIN(_12404_),
    .COUT(_12405_),
    .SUM(_12406_));
 sky130_fd_sc_hd__fa_1 _27383_ (.A(\hash.CA1.k_i2[9] ),
    .B(\hash.CA1.w_i2[9] ),
    .CIN(_12407_),
    .COUT(_12408_),
    .SUM(_12409_));
 sky130_fd_sc_hd__fa_1 _27384_ (.A(\hash.CA1.k_i2[10] ),
    .B(\hash.CA1.w_i2[10] ),
    .CIN(_12410_),
    .COUT(_12411_),
    .SUM(_12412_));
 sky130_fd_sc_hd__fa_1 _27385_ (.A(_12413_),
    .B(_12414_),
    .CIN(_12415_),
    .COUT(_12416_),
    .SUM(_12417_));
 sky130_fd_sc_hd__fa_1 _27386_ (.A(_12418_),
    .B(_12419_),
    .CIN(_12420_),
    .COUT(_12421_),
    .SUM(_12422_));
 sky130_fd_sc_hd__fa_1 _27387_ (.A(\hash.CA1.k_i2[13] ),
    .B(\hash.CA1.w_i2[13] ),
    .CIN(_12423_),
    .COUT(_12424_),
    .SUM(_12425_));
 sky130_fd_sc_hd__fa_1 _27388_ (.A(_12426_),
    .B(_12427_),
    .CIN(_12428_),
    .COUT(_12429_),
    .SUM(_12430_));
 sky130_fd_sc_hd__fa_1 _27389_ (.A(_12431_),
    .B(_12432_),
    .CIN(_12433_),
    .COUT(_12434_),
    .SUM(_12435_));
 sky130_fd_sc_hd__fa_1 _27390_ (.A(_12436_),
    .B(_12437_),
    .CIN(_12438_),
    .COUT(_12439_),
    .SUM(_12440_));
 sky130_fd_sc_hd__fa_1 _27391_ (.A(_12441_),
    .B(_12442_),
    .CIN(_12443_),
    .COUT(_12444_),
    .SUM(_12445_));
 sky130_fd_sc_hd__fa_1 _27392_ (.A(\hash.CA1.k_i2[18] ),
    .B(\hash.CA1.w_i2[18] ),
    .CIN(_12446_),
    .COUT(_12447_),
    .SUM(_12448_));
 sky130_fd_sc_hd__fa_1 _27393_ (.A(\hash.CA1.k_i2[19] ),
    .B(\hash.CA1.w_i2[19] ),
    .CIN(_12449_),
    .COUT(_12450_),
    .SUM(_12451_));
 sky130_fd_sc_hd__fa_1 _27394_ (.A(\hash.CA1.k_i2[20] ),
    .B(\hash.CA1.w_i2[20] ),
    .CIN(_12452_),
    .COUT(_12453_),
    .SUM(_12454_));
 sky130_fd_sc_hd__fa_1 _27395_ (.A(\hash.CA1.k_i2[21] ),
    .B(\hash.CA1.w_i2[21] ),
    .CIN(_12455_),
    .COUT(_12456_),
    .SUM(_12457_));
 sky130_fd_sc_hd__fa_1 _27396_ (.A(\hash.CA1.k_i2[22] ),
    .B(\hash.CA1.w_i2[22] ),
    .CIN(_12458_),
    .COUT(_12459_),
    .SUM(_12460_));
 sky130_fd_sc_hd__fa_1 _27397_ (.A(_12461_),
    .B(_12462_),
    .CIN(_12463_),
    .COUT(_12464_),
    .SUM(_12465_));
 sky130_fd_sc_hd__fa_1 _27398_ (.A(_12466_),
    .B(_12467_),
    .CIN(_12468_),
    .COUT(_12469_),
    .SUM(_12470_));
 sky130_fd_sc_hd__fa_1 _27399_ (.A(_12471_),
    .B(_12472_),
    .CIN(_12473_),
    .COUT(_12474_),
    .SUM(_12475_));
 sky130_fd_sc_hd__fa_1 _27400_ (.A(_12476_),
    .B(_12477_),
    .CIN(_12478_),
    .COUT(_12479_),
    .SUM(_12480_));
 sky130_fd_sc_hd__fa_1 _27401_ (.A(_12481_),
    .B(_12482_),
    .CIN(_12483_),
    .COUT(_12484_),
    .SUM(_12485_));
 sky130_fd_sc_hd__fa_1 _27402_ (.A(_12486_),
    .B(_12487_),
    .CIN(_12488_),
    .COUT(_12489_),
    .SUM(_12490_));
 sky130_fd_sc_hd__fa_1 _27403_ (.A(\hash.CA1.k_i2[29] ),
    .B(\hash.CA1.w_i2[29] ),
    .CIN(_12491_),
    .COUT(_12492_),
    .SUM(_12493_));
 sky130_fd_sc_hd__fa_1 _27404_ (.A(\hash.CA1.k_i2[30] ),
    .B(\hash.CA1.w_i2[30] ),
    .CIN(_12494_),
    .COUT(_12495_),
    .SUM(_12496_));
 sky130_fd_sc_hd__fa_4 _27405_ (.A(\hash.CA1.k_i1[1] ),
    .B(\hash.CA1.w_i1[1] ),
    .CIN(_12497_),
    .COUT(_12498_),
    .SUM(_12499_));
 sky130_fd_sc_hd__fa_2 _27406_ (.A(_12502_),
    .B(_12501_),
    .CIN(_12500_),
    .COUT(_12503_),
    .SUM(_12504_));
 sky130_fd_sc_hd__fa_1 _27407_ (.A(_12504_),
    .B(_12499_),
    .CIN(_12505_),
    .COUT(_12506_),
    .SUM(_12507_));
 sky130_fd_sc_hd__fa_1 _27408_ (.A(_12508_),
    .B(_12509_),
    .CIN(_12510_),
    .COUT(_12511_),
    .SUM(_12512_));
 sky130_fd_sc_hd__fa_1 _27409_ (.A(_12513_),
    .B(_12514_),
    .CIN(_12515_),
    .COUT(_12516_),
    .SUM(_12517_));
 sky130_fd_sc_hd__fa_1 _27410_ (.A(_12518_),
    .B(_12519_),
    .CIN(_12520_),
    .COUT(_12521_),
    .SUM(_12522_));
 sky130_fd_sc_hd__fa_1 _27411_ (.A(_12523_),
    .B(_12524_),
    .CIN(_12525_),
    .COUT(_12526_),
    .SUM(_12527_));
 sky130_fd_sc_hd__fa_1 _27412_ (.A(_12528_),
    .B(_12529_),
    .CIN(_12530_),
    .COUT(_12531_),
    .SUM(_12532_));
 sky130_fd_sc_hd__fa_1 _27413_ (.A(_12533_),
    .B(_12534_),
    .CIN(_12535_),
    .COUT(_12536_),
    .SUM(_12537_));
 sky130_fd_sc_hd__fa_1 _27414_ (.A(_12538_),
    .B(_12539_),
    .CIN(_12540_),
    .COUT(_12541_),
    .SUM(_12542_));
 sky130_fd_sc_hd__fa_2 _27415_ (.A(_12545_),
    .B(_12544_),
    .CIN(_12543_),
    .COUT(_12546_),
    .SUM(_12547_));
 sky130_fd_sc_hd__fa_1 _27416_ (.A(_12550_),
    .B(_12549_),
    .CIN(_12548_),
    .COUT(_12551_),
    .SUM(_12552_));
 sky130_fd_sc_hd__fa_1 _27417_ (.A(_12553_),
    .B(_12554_),
    .CIN(_12555_),
    .COUT(_12556_),
    .SUM(_12557_));
 sky130_fd_sc_hd__fa_1 _27418_ (.A(_12560_),
    .B(_12559_),
    .CIN(_12558_),
    .COUT(_12561_),
    .SUM(_12562_));
 sky130_fd_sc_hd__fa_1 _27419_ (.A(_12563_),
    .B(_12564_),
    .CIN(_12565_),
    .COUT(_12566_),
    .SUM(_12567_));
 sky130_fd_sc_hd__fa_1 _27420_ (.A(_12570_),
    .B(_12569_),
    .CIN(_12568_),
    .COUT(_12571_),
    .SUM(_12572_));
 sky130_fd_sc_hd__fa_1 _27421_ (.A(_12573_),
    .B(_12574_),
    .CIN(_12575_),
    .COUT(_12576_),
    .SUM(_12577_));
 sky130_fd_sc_hd__fa_1 _27422_ (.A(_12578_),
    .B(_12579_),
    .CIN(_12580_),
    .COUT(_12581_),
    .SUM(_12582_));
 sky130_fd_sc_hd__fa_1 _27423_ (.A(_12583_),
    .B(_12584_),
    .CIN(_12585_),
    .COUT(_12586_),
    .SUM(_12587_));
 sky130_fd_sc_hd__fa_1 _27424_ (.A(_12588_),
    .B(_12589_),
    .CIN(_06325_),
    .COUT(_12591_),
    .SUM(_12592_));
 sky130_fd_sc_hd__fa_1 _27425_ (.A(_12593_),
    .B(_12594_),
    .CIN(_12595_),
    .COUT(_12596_),
    .SUM(_12597_));
 sky130_fd_sc_hd__fa_1 _27426_ (.A(_12598_),
    .B(_12599_),
    .CIN(_12600_),
    .COUT(_12601_),
    .SUM(_12602_));
 sky130_fd_sc_hd__fa_1 _27427_ (.A(_12603_),
    .B(_12604_),
    .CIN(_12605_),
    .COUT(_12606_),
    .SUM(_12607_));
 sky130_fd_sc_hd__fa_1 _27428_ (.A(_12608_),
    .B(_12609_),
    .CIN(_12610_),
    .COUT(_12611_),
    .SUM(_12612_));
 sky130_fd_sc_hd__fa_1 _27429_ (.A(_12613_),
    .B(_12614_),
    .CIN(_12615_),
    .COUT(_12616_),
    .SUM(_12617_));
 sky130_fd_sc_hd__fa_1 _27430_ (.A(_12618_),
    .B(_12619_),
    .CIN(_12620_),
    .COUT(_12621_),
    .SUM(_12622_));
 sky130_fd_sc_hd__fa_1 _27431_ (.A(_12623_),
    .B(_12624_),
    .CIN(_12625_),
    .COUT(_12626_),
    .SUM(_12627_));
 sky130_fd_sc_hd__fa_1 _27432_ (.A(_12628_),
    .B(_12629_),
    .CIN(_12630_),
    .COUT(_12631_),
    .SUM(_12632_));
 sky130_fd_sc_hd__fa_1 _27433_ (.A(_12633_),
    .B(_12634_),
    .CIN(_12635_),
    .COUT(_12636_),
    .SUM(_12637_));
 sky130_fd_sc_hd__fa_1 _27434_ (.A(_12638_),
    .B(_12639_),
    .CIN(_12640_),
    .COUT(_12641_),
    .SUM(_12642_));
 sky130_fd_sc_hd__fa_1 _27435_ (.A(_12643_),
    .B(_12644_),
    .CIN(_12645_),
    .COUT(_12646_),
    .SUM(_12647_));
 sky130_fd_sc_hd__fa_1 _27436_ (.A(_12648_),
    .B(_12649_),
    .CIN(_12650_),
    .COUT(_12651_),
    .SUM(_12652_));
 sky130_fd_sc_hd__fa_1 _27437_ (.A(\hash.CA1.d[0] ),
    .B(_12653_),
    .CIN(_12654_),
    .COUT(_12655_),
    .SUM(_12656_));
 sky130_fd_sc_hd__fa_1 _27438_ (.A(_12657_),
    .B(_12499_),
    .CIN(_12505_),
    .COUT(_12658_),
    .SUM(_12659_));
 sky130_fd_sc_hd__fa_1 _27439_ (.A(_12660_),
    .B(_12661_),
    .CIN(_12662_),
    .COUT(_12663_),
    .SUM(_12664_));
 sky130_fd_sc_hd__fa_1 _27440_ (.A(_12665_),
    .B(_12666_),
    .CIN(_12667_),
    .COUT(_12668_),
    .SUM(_12669_));
 sky130_fd_sc_hd__fa_1 _27441_ (.A(_12670_),
    .B(_12669_),
    .CIN(_12671_),
    .COUT(_12672_),
    .SUM(_12673_));
 sky130_fd_sc_hd__fa_1 _27442_ (.A(_12514_),
    .B(_12674_),
    .CIN(_12515_),
    .COUT(_12675_),
    .SUM(_12676_));
 sky130_fd_sc_hd__fa_1 _27443_ (.A(_12668_),
    .B(_12676_),
    .CIN(_12513_),
    .COUT(_12677_),
    .SUM(_12678_));
 sky130_fd_sc_hd__fa_1 _27444_ (.A(_12519_),
    .B(_12679_),
    .CIN(_12520_),
    .COUT(_12680_),
    .SUM(_12681_));
 sky130_fd_sc_hd__fa_1 _27445_ (.A(_12675_),
    .B(_12681_),
    .CIN(_12518_),
    .COUT(_12682_),
    .SUM(_12683_));
 sky130_fd_sc_hd__fa_1 _27446_ (.A(_12524_),
    .B(_12684_),
    .CIN(_12525_),
    .COUT(_12685_),
    .SUM(_12686_));
 sky130_fd_sc_hd__fa_1 _27447_ (.A(_12680_),
    .B(_12687_),
    .CIN(_12688_),
    .COUT(_12689_),
    .SUM(_12690_));
 sky130_fd_sc_hd__fa_1 _27448_ (.A(_12691_),
    .B(_12692_),
    .CIN(_12693_),
    .COUT(_12694_),
    .SUM(_12695_));
 sky130_fd_sc_hd__fa_1 _27449_ (.A(_12696_),
    .B(_12695_),
    .CIN(_12697_),
    .COUT(_12698_),
    .SUM(_12699_));
 sky130_fd_sc_hd__fa_1 _27450_ (.A(_12700_),
    .B(_12701_),
    .CIN(_12702_),
    .COUT(_12703_),
    .SUM(_12704_));
 sky130_fd_sc_hd__fa_1 _27451_ (.A(_12694_),
    .B(_12704_),
    .CIN(_12705_),
    .COUT(_12706_),
    .SUM(_12707_));
 sky130_fd_sc_hd__fa_1 _27452_ (.A(_12539_),
    .B(_12708_),
    .CIN(_12540_),
    .COUT(_12709_),
    .SUM(_12710_));
 sky130_fd_sc_hd__fa_1 _27453_ (.A(_12703_),
    .B(_12710_),
    .CIN(_12538_),
    .COUT(_12711_),
    .SUM(_12712_));
 sky130_fd_sc_hd__fa_1 _27454_ (.A(_12713_),
    .B(_12714_),
    .CIN(_12715_),
    .COUT(_12716_),
    .SUM(_12717_));
 sky130_fd_sc_hd__fa_1 _27455_ (.A(_12718_),
    .B(_12719_),
    .CIN(_12720_),
    .COUT(_12721_),
    .SUM(_12722_));
 sky130_fd_sc_hd__fa_1 _27456_ (.A(_12549_),
    .B(_12723_),
    .CIN(_12550_),
    .COUT(_12724_),
    .SUM(_12725_));
 sky130_fd_sc_hd__fa_1 _27457_ (.A(_12726_),
    .B(_12727_),
    .CIN(net1098),
    .COUT(_12729_),
    .SUM(_12730_));
 sky130_fd_sc_hd__fa_1 _27458_ (.A(_12731_),
    .B(_12732_),
    .CIN(_12733_),
    .COUT(_12734_),
    .SUM(_12735_));
 sky130_fd_sc_hd__fa_1 _27459_ (.A(_12736_),
    .B(_12735_),
    .CIN(_12737_),
    .COUT(_12738_),
    .SUM(_12739_));
 sky130_fd_sc_hd__fa_1 _27460_ (.A(_12559_),
    .B(_06747_),
    .CIN(_12560_),
    .COUT(_12741_),
    .SUM(_12742_));
 sky130_fd_sc_hd__fa_1 _27461_ (.A(_12734_),
    .B(_12742_),
    .CIN(_12743_),
    .COUT(_12744_),
    .SUM(_12745_));
 sky130_fd_sc_hd__fa_1 _27462_ (.A(_12564_),
    .B(_12746_),
    .CIN(_12565_),
    .COUT(_12747_),
    .SUM(_12748_));
 sky130_fd_sc_hd__fa_1 _27463_ (.A(_12741_),
    .B(_12748_),
    .CIN(_12749_),
    .COUT(_12750_),
    .SUM(_12751_));
 sky130_fd_sc_hd__fa_1 _27464_ (.A(_12569_),
    .B(_12752_),
    .CIN(_12570_),
    .COUT(_12753_),
    .SUM(_12754_));
 sky130_fd_sc_hd__fa_1 _27465_ (.A(_12747_),
    .B(_12755_),
    .CIN(_12756_),
    .COUT(_12757_),
    .SUM(_12758_));
 sky130_fd_sc_hd__fa_1 _27466_ (.A(_12574_),
    .B(_12759_),
    .CIN(_12575_),
    .COUT(_12760_),
    .SUM(_12761_));
 sky130_fd_sc_hd__fa_1 _27467_ (.A(_12762_),
    .B(_12763_),
    .CIN(_12764_),
    .COUT(_12765_),
    .SUM(_12766_));
 sky130_fd_sc_hd__fa_1 _27468_ (.A(_12579_),
    .B(_12767_),
    .CIN(_12580_),
    .COUT(_12768_),
    .SUM(_12769_));
 sky130_fd_sc_hd__fa_1 _27469_ (.A(_12770_),
    .B(_12769_),
    .CIN(_12771_),
    .COUT(_12772_),
    .SUM(_12773_));
 sky130_fd_sc_hd__fa_1 _27470_ (.A(_12584_),
    .B(_12774_),
    .CIN(_12585_),
    .COUT(_12775_),
    .SUM(_12776_));
 sky130_fd_sc_hd__fa_1 _27471_ (.A(_12768_),
    .B(_12776_),
    .CIN(_12777_),
    .COUT(_12778_),
    .SUM(_12779_));
 sky130_fd_sc_hd__fa_1 _27472_ (.A(_12589_),
    .B(_12780_),
    .CIN(_06325_),
    .COUT(_12781_),
    .SUM(_12782_));
 sky130_fd_sc_hd__fa_1 _27473_ (.A(_12775_),
    .B(_12782_),
    .CIN(_12783_),
    .COUT(_12784_),
    .SUM(_12785_));
 sky130_fd_sc_hd__fa_1 _27474_ (.A(_12594_),
    .B(_12786_),
    .CIN(_12595_),
    .COUT(_12787_),
    .SUM(_12788_));
 sky130_fd_sc_hd__fa_1 _27475_ (.A(_12781_),
    .B(_12788_),
    .CIN(_12789_),
    .COUT(_12790_),
    .SUM(_12791_));
 sky130_fd_sc_hd__fa_1 _27476_ (.A(_12792_),
    .B(_12793_),
    .CIN(_12794_),
    .COUT(_12795_),
    .SUM(_12796_));
 sky130_fd_sc_hd__fa_1 _27477_ (.A(_12787_),
    .B(_12797_),
    .CIN(_12798_),
    .COUT(_12799_),
    .SUM(_12800_));
 sky130_fd_sc_hd__fa_1 _27478_ (.A(_12801_),
    .B(_12802_),
    .CIN(_12803_),
    .COUT(_12804_),
    .SUM(_12805_));
 sky130_fd_sc_hd__fa_1 _27479_ (.A(_12806_),
    .B(_12805_),
    .CIN(_12807_),
    .COUT(_12808_),
    .SUM(_12809_));
 sky130_fd_sc_hd__fa_1 _27480_ (.A(_12609_),
    .B(_12810_),
    .CIN(_12610_),
    .COUT(_12811_),
    .SUM(_12812_));
 sky130_fd_sc_hd__fa_1 _27481_ (.A(_12804_),
    .B(_12813_),
    .CIN(_12814_),
    .COUT(_12815_),
    .SUM(_12816_));
 sky130_fd_sc_hd__fa_1 _27482_ (.A(_12817_),
    .B(_12818_),
    .CIN(_12819_),
    .COUT(_12820_),
    .SUM(_12821_));
 sky130_fd_sc_hd__fa_1 _27483_ (.A(_12822_),
    .B(_12821_),
    .CIN(_12823_),
    .COUT(_12824_),
    .SUM(_12825_));
 sky130_fd_sc_hd__fa_1 _27484_ (.A(_12619_),
    .B(_12826_),
    .CIN(_12620_),
    .COUT(_12827_),
    .SUM(_12828_));
 sky130_fd_sc_hd__fa_1 _27485_ (.A(_12820_),
    .B(_12830_),
    .CIN(_12829_),
    .COUT(_12831_),
    .SUM(_12832_));
 sky130_fd_sc_hd__fa_1 _27486_ (.A(_12833_),
    .B(_12834_),
    .CIN(_12835_),
    .COUT(_12836_),
    .SUM(_12837_));
 sky130_fd_sc_hd__fa_1 _27487_ (.A(_12838_),
    .B(_12837_),
    .CIN(_12839_),
    .COUT(_12840_),
    .SUM(_12841_));
 sky130_fd_sc_hd__fa_1 _27488_ (.A(_12629_),
    .B(_12842_),
    .CIN(_12630_),
    .COUT(_12843_),
    .SUM(_12844_));
 sky130_fd_sc_hd__fa_1 _27489_ (.A(_12836_),
    .B(_12844_),
    .CIN(_12845_),
    .COUT(_12846_),
    .SUM(_12847_));
 sky130_fd_sc_hd__fa_1 _27490_ (.A(_12848_),
    .B(_12849_),
    .CIN(_12850_),
    .COUT(_12851_),
    .SUM(_12852_));
 sky130_fd_sc_hd__fa_1 _27491_ (.A(_12843_),
    .B(_12852_),
    .CIN(_12853_),
    .COUT(_12854_),
    .SUM(_12855_));
 sky130_fd_sc_hd__fa_1 _27492_ (.A(_12856_),
    .B(_12857_),
    .CIN(_12858_),
    .COUT(_12859_),
    .SUM(_12860_));
 sky130_fd_sc_hd__fa_1 _27493_ (.A(_12851_),
    .B(_12860_),
    .CIN(_12861_),
    .COUT(_12862_),
    .SUM(_12863_));
 sky130_fd_sc_hd__fa_1 _27494_ (.A(_12644_),
    .B(_12864_),
    .CIN(_12645_),
    .COUT(_12865_),
    .SUM(_12866_));
 sky130_fd_sc_hd__fa_1 _27495_ (.A(_12859_),
    .B(_12866_),
    .CIN(_12867_),
    .COUT(_12868_),
    .SUM(_12869_));
 sky130_fd_sc_hd__fa_1 _27496_ (.A(_12870_),
    .B(_12871_),
    .CIN(_12872_),
    .COUT(_12873_),
    .SUM(_12874_));
 sky130_fd_sc_hd__fa_1 _27497_ (.A(_12875_),
    .B(_12876_),
    .CIN(_12648_),
    .COUT(_12877_),
    .SUM(_12878_));
 sky130_fd_sc_hd__fa_1 _27498_ (.A(_12879_),
    .B(_12880_),
    .CIN(_12881_),
    .COUT(_12882_),
    .SUM(_12883_));
 sky130_fd_sc_hd__fa_1 _27499_ (.A(_12884_),
    .B(_12663_),
    .CIN(_12673_),
    .COUT(_12885_),
    .SUM(_12886_));
 sky130_fd_sc_hd__fa_1 _27500_ (.A(_12653_),
    .B(_12887_),
    .CIN(_12654_),
    .COUT(_12888_),
    .SUM(\hash.CA1.p3[0] ));
 sky130_fd_sc_hd__fa_1 _27501_ (.A(_12889_),
    .B(_12890_),
    .CIN(_12891_),
    .COUT(_12892_),
    .SUM(_12893_));
 sky130_fd_sc_hd__fa_1 _27502_ (.A(_00721_),
    .B(_12894_),
    .CIN(_12895_),
    .COUT(_12896_),
    .SUM(_12897_));
 sky130_fd_sc_hd__ha_4 _27503_ (.A(_00656_),
    .B(_12900_),
    .COUT(_12901_),
    .SUM(_00657_));
 sky130_fd_sc_hd__ha_4 _27504_ (.A(_00656_),
    .B(\count_hash2[2] ),
    .COUT(_12902_),
    .SUM(_12903_));
 sky130_fd_sc_hd__ha_4 _27505_ (.A(\count_hash2[1] ),
    .B(_12900_),
    .COUT(_12904_),
    .SUM(_12905_));
 sky130_fd_sc_hd__ha_4 _27506_ (.A(\count_hash2[1] ),
    .B(\count_hash2[2] ),
    .COUT(_12906_),
    .SUM(_12907_));
 sky130_fd_sc_hd__ha_4 _27507_ (.A(\count_hash2[1] ),
    .B(\count_hash2[2] ),
    .COUT(_12908_),
    .SUM(_12909_));
 sky130_fd_sc_hd__ha_4 _27508_ (.A(_00654_),
    .B(_12910_),
    .COUT(_12911_),
    .SUM(_00655_));
 sky130_fd_sc_hd__ha_4 _27509_ (.A(_00654_),
    .B(\count_hash1[2] ),
    .COUT(_12912_),
    .SUM(_12913_));
 sky130_fd_sc_hd__ha_1 _27510_ (.A(_00654_),
    .B(\count_hash1[2] ),
    .COUT(_12914_),
    .SUM(_12915_));
 sky130_fd_sc_hd__ha_4 _27511_ (.A(net371),
    .B(_12910_),
    .COUT(_12916_),
    .SUM(_12917_));
 sky130_fd_sc_hd__ha_4 _27512_ (.A(net371),
    .B(\count_hash1[2] ),
    .COUT(_12918_),
    .SUM(_12919_));
 sky130_fd_sc_hd__ha_4 _27513_ (.A(\count_hash1[1] ),
    .B(\count_hash1[2] ),
    .COUT(_12920_),
    .SUM(_12921_));
 sky130_fd_sc_hd__ha_4 _27514_ (.A(\hash.CA2.p3[0] ),
    .B(\hash.CA2.p1[0] ),
    .COUT(_12080_),
    .SUM(_12922_));
 sky130_fd_sc_hd__ha_4 _27515_ (.A(\hash.CA2.p1[2] ),
    .B(\hash.CA2.p3[2] ),
    .COUT(_12923_),
    .SUM(_12924_));
 sky130_fd_sc_hd__ha_1 _27516_ (.A(\hash.CA2.p1[1] ),
    .B(\hash.CA2.p3[1] ),
    .COUT(_12925_),
    .SUM(_12926_));
 sky130_fd_sc_hd__ha_4 _27517_ (.A(\hash.CA2.p1[7] ),
    .B(\hash.CA2.p3[7] ),
    .COUT(_12927_),
    .SUM(_12928_));
 sky130_fd_sc_hd__ha_2 _27518_ (.A(\hash.CA2.p1[6] ),
    .B(\hash.CA2.p3[6] ),
    .COUT(_12929_),
    .SUM(_12930_));
 sky130_fd_sc_hd__ha_2 _27519_ (.A(\hash.CA2.p1[5] ),
    .B(\hash.CA2.p3[5] ),
    .COUT(_12931_),
    .SUM(_12932_));
 sky130_fd_sc_hd__ha_2 _27520_ (.A(\hash.CA2.p1[4] ),
    .B(\hash.CA2.p3[4] ),
    .COUT(_12933_),
    .SUM(_12934_));
 sky130_fd_sc_hd__ha_4 _27521_ (.A(\hash.CA2.p1[3] ),
    .B(\hash.CA2.p3[3] ),
    .COUT(_12935_),
    .SUM(_12936_));
 sky130_fd_sc_hd__ha_4 _27522_ (.A(\hash.CA2.p1[9] ),
    .B(\hash.CA2.p3[9] ),
    .COUT(_12937_),
    .SUM(_12938_));
 sky130_fd_sc_hd__ha_4 _27523_ (.A(\hash.CA2.p1[8] ),
    .B(\hash.CA2.p3[8] ),
    .COUT(_12939_),
    .SUM(_12940_));
 sky130_fd_sc_hd__ha_1 _27524_ (.A(\hash.CA2.p1[10] ),
    .B(\hash.CA2.p3[10] ),
    .COUT(_12941_),
    .SUM(_12942_));
 sky130_fd_sc_hd__ha_4 _27525_ (.A(\hash.CA2.p1[11] ),
    .B(\hash.CA2.p3[11] ),
    .COUT(_12943_),
    .SUM(_12944_));
 sky130_fd_sc_hd__ha_2 _27526_ (.A(\hash.CA2.p1[13] ),
    .B(\hash.CA2.p3[13] ),
    .COUT(_12945_),
    .SUM(_12946_));
 sky130_fd_sc_hd__ha_4 _27527_ (.A(\hash.CA2.p1[12] ),
    .B(\hash.CA2.p3[12] ),
    .COUT(_12947_),
    .SUM(_12948_));
 sky130_fd_sc_hd__ha_1 _27528_ (.A(\hash.CA2.p1[15] ),
    .B(\hash.CA2.p3[15] ),
    .COUT(_12949_),
    .SUM(_12950_));
 sky130_fd_sc_hd__ha_1 _27529_ (.A(\hash.CA2.p1[14] ),
    .B(\hash.CA2.p3[14] ),
    .COUT(_12951_),
    .SUM(_12952_));
 sky130_fd_sc_hd__ha_4 _27530_ (.A(\hash.CA2.p1[16] ),
    .B(\hash.CA2.p3[16] ),
    .COUT(_12953_),
    .SUM(_12954_));
 sky130_fd_sc_hd__ha_2 _27531_ (.A(\hash.CA2.p1[17] ),
    .B(\hash.CA2.p3[17] ),
    .COUT(_12955_),
    .SUM(_12956_));
 sky130_fd_sc_hd__ha_1 _27532_ (.A(\hash.CA2.p1[18] ),
    .B(\hash.CA2.p3[18] ),
    .COUT(_12957_),
    .SUM(_12958_));
 sky130_fd_sc_hd__ha_4 _27533_ (.A(\hash.CA2.p1[21] ),
    .B(\hash.CA2.p3[21] ),
    .COUT(_12959_),
    .SUM(_12960_));
 sky130_fd_sc_hd__ha_4 _27534_ (.A(\hash.CA2.p1[20] ),
    .B(\hash.CA2.p3[20] ),
    .COUT(_12961_),
    .SUM(_12962_));
 sky130_fd_sc_hd__ha_4 _27535_ (.A(\hash.CA2.p1[19] ),
    .B(\hash.CA2.p3[19] ),
    .COUT(_12963_),
    .SUM(_12964_));
 sky130_fd_sc_hd__ha_4 _27536_ (.A(\hash.CA2.p1[22] ),
    .B(\hash.CA2.p3[22] ),
    .COUT(_12965_),
    .SUM(_12966_));
 sky130_fd_sc_hd__ha_4 _27537_ (.A(\hash.CA2.p1[24] ),
    .B(\hash.CA2.p3[24] ),
    .COUT(_12967_),
    .SUM(_12968_));
 sky130_fd_sc_hd__ha_4 _27538_ (.A(\hash.CA2.p1[23] ),
    .B(\hash.CA2.p3[23] ),
    .COUT(_12969_),
    .SUM(_12970_));
 sky130_fd_sc_hd__ha_4 _27539_ (.A(\hash.CA2.p1[25] ),
    .B(\hash.CA2.p3[25] ),
    .COUT(_12971_),
    .SUM(_12972_));
 sky130_fd_sc_hd__ha_4 _27540_ (.A(\hash.CA2.p1[27] ),
    .B(\hash.CA2.p3[27] ),
    .COUT(_12973_),
    .SUM(_12974_));
 sky130_fd_sc_hd__ha_4 _27541_ (.A(\hash.CA2.p1[26] ),
    .B(\hash.CA2.p3[26] ),
    .COUT(_12975_),
    .SUM(_12976_));
 sky130_fd_sc_hd__ha_4 _27542_ (.A(\hash.CA2.p1[28] ),
    .B(\hash.CA2.p3[28] ),
    .COUT(_12977_),
    .SUM(_12978_));
 sky130_fd_sc_hd__ha_1 _27543_ (.A(\hash.CA2.p1[29] ),
    .B(\hash.CA2.p3[29] ),
    .COUT(_12979_),
    .SUM(_12980_));
 sky130_fd_sc_hd__ha_1 _27544_ (.A(\hash.CA2.p1[30] ),
    .B(\hash.CA2.p3[30] ),
    .COUT(_12981_),
    .SUM(_12982_));
 sky130_fd_sc_hd__ha_1 _27545_ (.A(_12983_),
    .B(_12984_),
    .COUT(_12985_),
    .SUM(_12986_));
 sky130_fd_sc_hd__ha_1 _27546_ (.A(_12985_),
    .B(_12987_),
    .COUT(_12988_),
    .SUM(_12989_));
 sky130_fd_sc_hd__ha_1 _27547_ (.A(_12990_),
    .B(_12991_),
    .COUT(_12992_),
    .SUM(_12993_));
 sky130_fd_sc_hd__ha_2 _27548_ (.A(_12994_),
    .B(_12995_),
    .COUT(_12996_),
    .SUM(_12997_));
 sky130_fd_sc_hd__ha_1 _27549_ (.A(_12998_),
    .B(_12999_),
    .COUT(_13000_),
    .SUM(_13001_));
 sky130_fd_sc_hd__ha_1 _27550_ (.A(_13002_),
    .B(_13003_),
    .COUT(_13004_),
    .SUM(_13005_));
 sky130_fd_sc_hd__ha_1 _27551_ (.A(_13006_),
    .B(_13007_),
    .COUT(_13008_),
    .SUM(_13009_));
 sky130_fd_sc_hd__ha_4 _27552_ (.A(_13010_),
    .B(_13011_),
    .COUT(_13012_),
    .SUM(_13013_));
 sky130_fd_sc_hd__ha_4 _27553_ (.A(_13014_),
    .B(_13015_),
    .COUT(_13016_),
    .SUM(_13017_));
 sky130_fd_sc_hd__ha_4 _27554_ (.A(_13018_),
    .B(_13019_),
    .COUT(_13020_),
    .SUM(_13021_));
 sky130_fd_sc_hd__ha_4 _27555_ (.A(_13022_),
    .B(_13023_),
    .COUT(_13024_),
    .SUM(_13025_));
 sky130_fd_sc_hd__ha_4 _27556_ (.A(_13026_),
    .B(_13027_),
    .COUT(_13028_),
    .SUM(_13029_));
 sky130_fd_sc_hd__ha_1 _27557_ (.A(_13030_),
    .B(_13031_),
    .COUT(_13032_),
    .SUM(_13033_));
 sky130_fd_sc_hd__ha_1 _27558_ (.A(_13034_),
    .B(_13035_),
    .COUT(_13036_),
    .SUM(_13037_));
 sky130_fd_sc_hd__ha_1 _27559_ (.A(_13038_),
    .B(_13039_),
    .COUT(_13040_),
    .SUM(_13041_));
 sky130_fd_sc_hd__ha_1 _27560_ (.A(_13042_),
    .B(_13043_),
    .COUT(_13044_),
    .SUM(_13045_));
 sky130_fd_sc_hd__ha_1 _27561_ (.A(_13046_),
    .B(_13047_),
    .COUT(_13048_),
    .SUM(_13049_));
 sky130_fd_sc_hd__ha_1 _27562_ (.A(_13050_),
    .B(_13051_),
    .COUT(_13052_),
    .SUM(_13053_));
 sky130_fd_sc_hd__ha_1 _27563_ (.A(_13054_),
    .B(_13055_),
    .COUT(_13056_),
    .SUM(_13057_));
 sky130_fd_sc_hd__ha_1 _27564_ (.A(_13058_),
    .B(_13059_),
    .COUT(_13060_),
    .SUM(_13061_));
 sky130_fd_sc_hd__ha_4 _27565_ (.A(_13062_),
    .B(_13063_),
    .COUT(_13064_),
    .SUM(_13065_));
 sky130_fd_sc_hd__ha_1 _27566_ (.A(_13066_),
    .B(_13067_),
    .COUT(_13068_),
    .SUM(_13069_));
 sky130_fd_sc_hd__ha_4 _27567_ (.A(_13070_),
    .B(_13071_),
    .COUT(_13072_),
    .SUM(_13073_));
 sky130_fd_sc_hd__ha_1 _27568_ (.A(_13074_),
    .B(_13075_),
    .COUT(_13076_),
    .SUM(_13077_));
 sky130_fd_sc_hd__ha_1 _27569_ (.A(_13078_),
    .B(_13079_),
    .COUT(_13080_),
    .SUM(_13081_));
 sky130_fd_sc_hd__ha_1 _27570_ (.A(_13082_),
    .B(_13083_),
    .COUT(_13084_),
    .SUM(_13085_));
 sky130_fd_sc_hd__ha_4 _27571_ (.A(_13086_),
    .B(_13087_),
    .COUT(_13088_),
    .SUM(_13089_));
 sky130_fd_sc_hd__ha_4 _27572_ (.A(_13090_),
    .B(_13091_),
    .COUT(_13092_),
    .SUM(_13093_));
 sky130_fd_sc_hd__ha_4 _27573_ (.A(_13094_),
    .B(_13095_),
    .COUT(_13096_),
    .SUM(_13097_));
 sky130_fd_sc_hd__ha_4 _27574_ (.A(_13098_),
    .B(_13099_),
    .COUT(_13100_),
    .SUM(_13101_));
 sky130_fd_sc_hd__ha_4 _27575_ (.A(_13102_),
    .B(_13103_),
    .COUT(_13104_),
    .SUM(_13105_));
 sky130_fd_sc_hd__ha_1 _27576_ (.A(_13106_),
    .B(_13107_),
    .COUT(_13108_),
    .SUM(_13109_));
 sky130_fd_sc_hd__ha_1 _27577_ (.A(_13108_),
    .B(_13110_),
    .COUT(_13111_),
    .SUM(_13112_));
 sky130_fd_sc_hd__ha_1 _27578_ (.A(_13113_),
    .B(_13114_),
    .COUT(_13115_),
    .SUM(_13116_));
 sky130_fd_sc_hd__ha_1 _27579_ (.A(_13117_),
    .B(_13118_),
    .COUT(_13119_),
    .SUM(_13120_));
 sky130_fd_sc_hd__ha_1 _27580_ (.A(_13121_),
    .B(_13122_),
    .COUT(_13123_),
    .SUM(_13124_));
 sky130_fd_sc_hd__ha_1 _27581_ (.A(_13125_),
    .B(_13126_),
    .COUT(_13127_),
    .SUM(_13128_));
 sky130_fd_sc_hd__ha_1 _27582_ (.A(_13129_),
    .B(_13130_),
    .COUT(_13131_),
    .SUM(_13132_));
 sky130_fd_sc_hd__ha_2 _27583_ (.A(_13133_),
    .B(_13134_),
    .COUT(_13135_),
    .SUM(_13136_));
 sky130_fd_sc_hd__ha_4 _27584_ (.A(_13137_),
    .B(_13138_),
    .COUT(_13139_),
    .SUM(_13140_));
 sky130_fd_sc_hd__ha_4 _27585_ (.A(_13141_),
    .B(_13142_),
    .COUT(_13143_),
    .SUM(_13144_));
 sky130_fd_sc_hd__ha_4 _27586_ (.A(_13145_),
    .B(_13146_),
    .COUT(_13147_),
    .SUM(_13148_));
 sky130_fd_sc_hd__ha_4 _27587_ (.A(_13149_),
    .B(_13150_),
    .COUT(_13151_),
    .SUM(_13152_));
 sky130_fd_sc_hd__ha_2 _27588_ (.A(_13153_),
    .B(_13154_),
    .COUT(_13155_),
    .SUM(_13156_));
 sky130_fd_sc_hd__ha_1 _27589_ (.A(_13157_),
    .B(_13158_),
    .COUT(_13159_),
    .SUM(_13160_));
 sky130_fd_sc_hd__ha_1 _27590_ (.A(_13161_),
    .B(_13162_),
    .COUT(_13163_),
    .SUM(_13164_));
 sky130_fd_sc_hd__ha_1 _27591_ (.A(_13165_),
    .B(_13166_),
    .COUT(_13167_),
    .SUM(_13168_));
 sky130_fd_sc_hd__ha_1 _27592_ (.A(_13169_),
    .B(_13170_),
    .COUT(_13171_),
    .SUM(_13172_));
 sky130_fd_sc_hd__ha_4 _27593_ (.A(_13173_),
    .B(_13174_),
    .COUT(_13175_),
    .SUM(_13176_));
 sky130_fd_sc_hd__ha_4 _27594_ (.A(_13177_),
    .B(_13178_),
    .COUT(_13179_),
    .SUM(_13180_));
 sky130_fd_sc_hd__ha_4 _27595_ (.A(_13181_),
    .B(_13182_),
    .COUT(_13183_),
    .SUM(_13184_));
 sky130_fd_sc_hd__ha_2 _27596_ (.A(_13185_),
    .B(_13186_),
    .COUT(_13187_),
    .SUM(_13188_));
 sky130_fd_sc_hd__ha_1 _27597_ (.A(_13189_),
    .B(_13190_),
    .COUT(_13191_),
    .SUM(_13192_));
 sky130_fd_sc_hd__ha_4 _27598_ (.A(_13193_),
    .B(_13194_),
    .COUT(_13195_),
    .SUM(_13196_));
 sky130_fd_sc_hd__ha_2 _27599_ (.A(_13197_),
    .B(_13198_),
    .COUT(_13199_),
    .SUM(_13200_));
 sky130_fd_sc_hd__ha_1 _27600_ (.A(_13201_),
    .B(_13202_),
    .COUT(_13203_),
    .SUM(_13204_));
 sky130_fd_sc_hd__ha_1 _27601_ (.A(_13205_),
    .B(_13206_),
    .COUT(_13207_),
    .SUM(_13208_));
 sky130_fd_sc_hd__ha_4 _27602_ (.A(_13209_),
    .B(_13210_),
    .COUT(_13211_),
    .SUM(_13212_));
 sky130_fd_sc_hd__ha_4 _27603_ (.A(_13213_),
    .B(_13214_),
    .COUT(_13215_),
    .SUM(_13216_));
 sky130_fd_sc_hd__ha_1 _27604_ (.A(_13217_),
    .B(_13218_),
    .COUT(_13219_),
    .SUM(_13220_));
 sky130_fd_sc_hd__ha_1 _27605_ (.A(_13221_),
    .B(_13222_),
    .COUT(_13223_),
    .SUM(_13224_));
 sky130_fd_sc_hd__ha_1 _27606_ (.A(_13225_),
    .B(_13226_),
    .COUT(_13227_),
    .SUM(_13228_));
 sky130_fd_sc_hd__ha_4 _27607_ (.A(_13230_),
    .B(_13229_),
    .COUT(_13231_),
    .SUM(_13232_));
 sky130_fd_sc_hd__ha_1 _27608_ (.A(\hash.CA2.p4[0] ),
    .B(_13233_),
    .COUT(_13234_),
    .SUM(_13235_));
 sky130_fd_sc_hd__ha_4 _27609_ (.A(_13236_),
    .B(_13237_),
    .COUT(_13238_),
    .SUM(_13239_));
 sky130_fd_sc_hd__ha_1 _27610_ (.A(_13234_),
    .B(_12095_),
    .COUT(_13240_),
    .SUM(_13241_));
 sky130_fd_sc_hd__ha_4 _27611_ (.A(_13243_),
    .B(_13242_),
    .COUT(_13244_),
    .SUM(_13245_));
 sky130_fd_sc_hd__ha_1 _27612_ (.A(_12094_),
    .B(_12104_),
    .COUT(_13247_),
    .SUM(_13248_));
 sky130_fd_sc_hd__ha_4 _27613_ (.A(_13249_),
    .B(_13250_),
    .COUT(_13251_),
    .SUM(_13252_));
 sky130_fd_sc_hd__ha_1 _27614_ (.A(_12103_),
    .B(_12118_),
    .COUT(_13254_),
    .SUM(_13255_));
 sky130_fd_sc_hd__ha_4 _27615_ (.A(_13256_),
    .B(_13257_),
    .COUT(_13258_),
    .SUM(_13259_));
 sky130_fd_sc_hd__ha_4 _27616_ (.A(_12117_),
    .B(_12127_),
    .COUT(_13261_),
    .SUM(_13262_));
 sky130_fd_sc_hd__ha_4 _27617_ (.A(_13263_),
    .B(_13264_),
    .COUT(_13265_),
    .SUM(_13266_));
 sky130_fd_sc_hd__ha_2 _27618_ (.A(_12126_),
    .B(_12136_),
    .COUT(_13268_),
    .SUM(_13269_));
 sky130_fd_sc_hd__ha_4 _27619_ (.A(_13270_),
    .B(_13271_),
    .COUT(_13272_),
    .SUM(_13273_));
 sky130_fd_sc_hd__ha_2 _27620_ (.A(_12135_),
    .B(_12145_),
    .COUT(_13275_),
    .SUM(_13276_));
 sky130_fd_sc_hd__ha_4 _27621_ (.A(_13277_),
    .B(_13278_),
    .COUT(_13279_),
    .SUM(_13280_));
 sky130_fd_sc_hd__ha_4 _27622_ (.A(_12144_),
    .B(_12154_),
    .COUT(_13282_),
    .SUM(_13283_));
 sky130_fd_sc_hd__ha_2 _27623_ (.A(_13284_),
    .B(_13285_),
    .COUT(_13286_),
    .SUM(_13287_));
 sky130_fd_sc_hd__ha_4 _27624_ (.A(_12153_),
    .B(_12163_),
    .COUT(_13289_),
    .SUM(_13290_));
 sky130_fd_sc_hd__ha_4 _27625_ (.A(_13291_),
    .B(_13292_),
    .COUT(_13293_),
    .SUM(_13294_));
 sky130_fd_sc_hd__ha_4 _27626_ (.A(_12162_),
    .B(_12172_),
    .COUT(_13296_),
    .SUM(_13297_));
 sky130_fd_sc_hd__ha_4 _27627_ (.A(_13298_),
    .B(_13299_),
    .COUT(_13300_),
    .SUM(_13301_));
 sky130_fd_sc_hd__ha_1 _27628_ (.A(_12171_),
    .B(_12181_),
    .COUT(_13303_),
    .SUM(_13304_));
 sky130_fd_sc_hd__ha_4 _27629_ (.A(_13305_),
    .B(_13306_),
    .COUT(_13307_),
    .SUM(_13308_));
 sky130_fd_sc_hd__ha_4 _27630_ (.A(_12180_),
    .B(_12190_),
    .COUT(_13310_),
    .SUM(_13311_));
 sky130_fd_sc_hd__ha_4 _27631_ (.A(_13312_),
    .B(_13313_),
    .COUT(_13314_),
    .SUM(_13315_));
 sky130_fd_sc_hd__ha_4 _27632_ (.A(_12189_),
    .B(_12199_),
    .COUT(_13317_),
    .SUM(_13318_));
 sky130_fd_sc_hd__ha_4 _27633_ (.A(_13319_),
    .B(_13320_),
    .COUT(_13321_),
    .SUM(_13322_));
 sky130_fd_sc_hd__ha_4 _27634_ (.A(_12198_),
    .B(_12208_),
    .COUT(_13324_),
    .SUM(_13325_));
 sky130_fd_sc_hd__ha_4 _27635_ (.A(_13326_),
    .B(_13327_),
    .COUT(_13328_),
    .SUM(_13329_));
 sky130_fd_sc_hd__ha_4 _27636_ (.A(_12207_),
    .B(_12217_),
    .COUT(_13331_),
    .SUM(_13332_));
 sky130_fd_sc_hd__ha_4 _27637_ (.A(_13333_),
    .B(_13334_),
    .COUT(_13335_),
    .SUM(_13336_));
 sky130_fd_sc_hd__ha_2 _27638_ (.A(_12216_),
    .B(_12226_),
    .COUT(_13338_),
    .SUM(_13339_));
 sky130_fd_sc_hd__ha_4 _27639_ (.A(_13340_),
    .B(_13341_),
    .COUT(_13342_),
    .SUM(_13343_));
 sky130_fd_sc_hd__ha_4 _27640_ (.A(_12225_),
    .B(_12235_),
    .COUT(_13345_),
    .SUM(_13346_));
 sky130_fd_sc_hd__ha_4 _27641_ (.A(_13347_),
    .B(_13348_),
    .COUT(_13349_),
    .SUM(_13350_));
 sky130_fd_sc_hd__ha_4 _27642_ (.A(_12234_),
    .B(_12244_),
    .COUT(_13352_),
    .SUM(_13353_));
 sky130_fd_sc_hd__ha_1 _27643_ (.A(_13354_),
    .B(_13355_),
    .COUT(_13356_),
    .SUM(_13357_));
 sky130_fd_sc_hd__ha_4 _27644_ (.A(_12243_),
    .B(_12253_),
    .COUT(_13359_),
    .SUM(_13360_));
 sky130_fd_sc_hd__ha_4 _27645_ (.A(_13361_),
    .B(_13362_),
    .COUT(_13363_),
    .SUM(_13364_));
 sky130_fd_sc_hd__ha_1 _27646_ (.A(_12252_),
    .B(_12262_),
    .COUT(_13366_),
    .SUM(_13367_));
 sky130_fd_sc_hd__ha_4 _27647_ (.A(_13368_),
    .B(_13369_),
    .COUT(_13370_),
    .SUM(_13371_));
 sky130_fd_sc_hd__ha_4 _27648_ (.A(_12261_),
    .B(_12271_),
    .COUT(_13373_),
    .SUM(_13374_));
 sky130_fd_sc_hd__ha_4 _27649_ (.A(_13375_),
    .B(_13376_),
    .COUT(_13377_),
    .SUM(_13378_));
 sky130_fd_sc_hd__ha_4 _27650_ (.A(_12270_),
    .B(_12280_),
    .COUT(_13380_),
    .SUM(_13381_));
 sky130_fd_sc_hd__ha_4 _27651_ (.A(_13382_),
    .B(_13383_),
    .COUT(_13384_),
    .SUM(_13385_));
 sky130_fd_sc_hd__ha_4 _27652_ (.A(_12279_),
    .B(_12289_),
    .COUT(_13387_),
    .SUM(_13388_));
 sky130_fd_sc_hd__ha_4 _27653_ (.A(_13389_),
    .B(_13390_),
    .COUT(_13391_),
    .SUM(_13392_));
 sky130_fd_sc_hd__ha_4 _27654_ (.A(_12288_),
    .B(_12298_),
    .COUT(_13394_),
    .SUM(_13395_));
 sky130_fd_sc_hd__ha_1 _27655_ (.A(_13396_),
    .B(_13397_),
    .COUT(_13398_),
    .SUM(_13399_));
 sky130_fd_sc_hd__ha_4 _27656_ (.A(_12297_),
    .B(_12307_),
    .COUT(_13401_),
    .SUM(_13402_));
 sky130_fd_sc_hd__ha_4 _27657_ (.A(_13403_),
    .B(_13404_),
    .COUT(_13405_),
    .SUM(_13406_));
 sky130_fd_sc_hd__ha_1 _27658_ (.A(_12306_),
    .B(_12316_),
    .COUT(_13408_),
    .SUM(_13409_));
 sky130_fd_sc_hd__ha_4 _27659_ (.A(_13410_),
    .B(_13411_),
    .COUT(_13412_),
    .SUM(_13413_));
 sky130_fd_sc_hd__ha_4 _27660_ (.A(_12315_),
    .B(_12325_),
    .COUT(_13415_),
    .SUM(_13416_));
 sky130_fd_sc_hd__ha_2 _27661_ (.A(_13417_),
    .B(_13418_),
    .COUT(_13419_),
    .SUM(_13420_));
 sky130_fd_sc_hd__ha_4 _27662_ (.A(_12324_),
    .B(_12334_),
    .COUT(_13422_),
    .SUM(_13423_));
 sky130_fd_sc_hd__ha_1 _27663_ (.A(_13424_),
    .B(_13425_),
    .COUT(_13426_),
    .SUM(_13427_));
 sky130_fd_sc_hd__ha_1 _27664_ (.A(_12333_),
    .B(_12343_),
    .COUT(_13429_),
    .SUM(_13430_));
 sky130_fd_sc_hd__ha_1 _27665_ (.A(_13431_),
    .B(_13432_),
    .COUT(_13433_),
    .SUM(_13434_));
 sky130_fd_sc_hd__ha_4 _27666_ (.A(_12342_),
    .B(_12352_),
    .COUT(_13436_),
    .SUM(_13437_));
 sky130_fd_sc_hd__ha_1 _27667_ (.A(_13438_),
    .B(_13439_),
    .COUT(_13440_),
    .SUM(_13441_));
 sky130_fd_sc_hd__ha_4 _27668_ (.A(_12351_),
    .B(_12361_),
    .COUT(_13443_),
    .SUM(_13444_));
 sky130_fd_sc_hd__ha_4 _27669_ (.A(\hash.CA2.p5[0] ),
    .B(_13232_),
    .COUT(_12362_),
    .SUM(_13445_));
 sky130_fd_sc_hd__ha_1 _27670_ (.A(\hash.CA2.p5[1] ),
    .B(_12363_),
    .COUT(_13446_),
    .SUM(_13447_));
 sky130_fd_sc_hd__ha_4 _27671_ (.A(\hash.CA2.p5[2] ),
    .B(_13246_),
    .COUT(_13448_),
    .SUM(_13449_));
 sky130_fd_sc_hd__ha_4 _27672_ (.A(\hash.CA2.p5[3] ),
    .B(_13253_),
    .COUT(_13450_),
    .SUM(_13451_));
 sky130_fd_sc_hd__ha_4 _27673_ (.A(\hash.CA2.p5[4] ),
    .B(_13260_),
    .COUT(_13452_),
    .SUM(_13453_));
 sky130_fd_sc_hd__ha_4 _27674_ (.A(\hash.CA2.p5[5] ),
    .B(_13267_),
    .COUT(_13454_),
    .SUM(_13455_));
 sky130_fd_sc_hd__ha_2 _27675_ (.A(\hash.CA2.p5[6] ),
    .B(_13274_),
    .COUT(_13456_),
    .SUM(_13457_));
 sky130_fd_sc_hd__ha_1 _27676_ (.A(\hash.CA2.p5[7] ),
    .B(_13281_),
    .COUT(_13458_),
    .SUM(_13459_));
 sky130_fd_sc_hd__ha_4 _27677_ (.A(_13288_),
    .B(\hash.CA2.p5[8] ),
    .COUT(_13460_),
    .SUM(_13461_));
 sky130_fd_sc_hd__ha_4 _27678_ (.A(\hash.CA2.p5[9] ),
    .B(_13295_),
    .COUT(_13462_),
    .SUM(_13463_));
 sky130_fd_sc_hd__ha_1 _27679_ (.A(\hash.CA2.p5[10] ),
    .B(_13302_),
    .COUT(_13464_),
    .SUM(_13465_));
 sky130_fd_sc_hd__ha_1 _27680_ (.A(\hash.CA2.p5[11] ),
    .B(_13309_),
    .COUT(_13466_),
    .SUM(_13467_));
 sky130_fd_sc_hd__ha_4 _27681_ (.A(\hash.CA2.p5[12] ),
    .B(_13316_),
    .COUT(_13468_),
    .SUM(_13469_));
 sky130_fd_sc_hd__ha_1 _27682_ (.A(\hash.CA2.p5[13] ),
    .B(_13323_),
    .COUT(_13470_),
    .SUM(_13471_));
 sky130_fd_sc_hd__ha_4 _27683_ (.A(\hash.CA2.p5[14] ),
    .B(_13330_),
    .COUT(_13472_),
    .SUM(_13473_));
 sky130_fd_sc_hd__ha_4 _27684_ (.A(\hash.CA2.p5[15] ),
    .B(_13337_),
    .COUT(_13474_),
    .SUM(_13475_));
 sky130_fd_sc_hd__ha_4 _27685_ (.A(\hash.CA2.p5[16] ),
    .B(_13344_),
    .COUT(_13476_),
    .SUM(_13477_));
 sky130_fd_sc_hd__ha_4 _27686_ (.A(\hash.CA2.p5[17] ),
    .B(_13351_),
    .COUT(_13478_),
    .SUM(_13479_));
 sky130_fd_sc_hd__ha_1 _27687_ (.A(\hash.CA2.p5[16] ),
    .B(_13344_),
    .COUT(_13480_),
    .SUM(_13481_));
 sky130_fd_sc_hd__ha_1 _27688_ (.A(\hash.CA2.p5[18] ),
    .B(_13358_),
    .COUT(_13482_),
    .SUM(_13483_));
 sky130_fd_sc_hd__ha_4 _27689_ (.A(\hash.CA2.p5[19] ),
    .B(_13365_),
    .COUT(_13484_),
    .SUM(_13485_));
 sky130_fd_sc_hd__ha_1 _27690_ (.A(\hash.CA2.p5[20] ),
    .B(_13372_),
    .COUT(_13486_),
    .SUM(_13487_));
 sky130_fd_sc_hd__ha_4 _27691_ (.A(\hash.CA2.p5[21] ),
    .B(_13379_),
    .COUT(_13488_),
    .SUM(_13489_));
 sky130_fd_sc_hd__ha_1 _27692_ (.A(\hash.CA2.p5[20] ),
    .B(_13372_),
    .COUT(_13490_),
    .SUM(_13491_));
 sky130_fd_sc_hd__ha_4 _27693_ (.A(_13386_),
    .B(\hash.CA2.p5[22] ),
    .COUT(_13492_),
    .SUM(_13493_));
 sky130_fd_sc_hd__ha_4 _27694_ (.A(\hash.CA2.p5[21] ),
    .B(net1068),
    .COUT(_13494_),
    .SUM(_13495_));
 sky130_fd_sc_hd__ha_4 _27695_ (.A(\hash.CA2.p5[23] ),
    .B(_13393_),
    .COUT(_13496_),
    .SUM(_13497_));
 sky130_fd_sc_hd__ha_4 _27696_ (.A(\hash.CA2.p5[22] ),
    .B(net1066),
    .COUT(_13498_),
    .SUM(_13499_));
 sky130_fd_sc_hd__ha_2 _27697_ (.A(\hash.CA2.p5[24] ),
    .B(_13400_),
    .COUT(_13500_),
    .SUM(_13501_));
 sky130_fd_sc_hd__ha_1 _27698_ (.A(\hash.CA2.p5[23] ),
    .B(_13393_),
    .COUT(_13502_),
    .SUM(_13503_));
 sky130_fd_sc_hd__ha_1 _27699_ (.A(\hash.CA2.p5[25] ),
    .B(_13407_),
    .COUT(_13504_),
    .SUM(_13505_));
 sky130_fd_sc_hd__ha_4 _27700_ (.A(_13414_),
    .B(\hash.CA2.p5[26] ),
    .COUT(_13506_),
    .SUM(_13507_));
 sky130_fd_sc_hd__ha_2 _27701_ (.A(\hash.CA2.p5[25] ),
    .B(_13407_),
    .COUT(_13508_),
    .SUM(_13509_));
 sky130_fd_sc_hd__ha_4 _27702_ (.A(\hash.CA2.p5[27] ),
    .B(_13421_),
    .COUT(_13510_),
    .SUM(_13511_));
 sky130_fd_sc_hd__ha_1 _27703_ (.A(\hash.CA2.p5[26] ),
    .B(_13414_),
    .COUT(_13512_),
    .SUM(_13513_));
 sky130_fd_sc_hd__ha_4 _27704_ (.A(\hash.CA2.p5[28] ),
    .B(_13428_),
    .COUT(_13514_),
    .SUM(_13515_));
 sky130_fd_sc_hd__ha_4 _27705_ (.A(\hash.CA2.p5[29] ),
    .B(_13435_),
    .COUT(_13516_),
    .SUM(_13517_));
 sky130_fd_sc_hd__ha_1 _27706_ (.A(\hash.CA2.p5[30] ),
    .B(_13442_),
    .COUT(_13518_),
    .SUM(_13519_));
 sky130_fd_sc_hd__ha_1 _27707_ (.A(net412),
    .B(net407),
    .COUT(_13520_),
    .SUM(_00643_));
 sky130_fd_sc_hd__ha_1 _27708_ (.A(net550),
    .B(\count15_1[2] ),
    .COUT(_13521_),
    .SUM(_00644_));
 sky130_fd_sc_hd__ha_1 _27709_ (.A(net490),
    .B(net485),
    .COUT(_13522_),
    .SUM(_00645_));
 sky130_fd_sc_hd__ha_1 _27710_ (.A(net430),
    .B(net541),
    .COUT(_13523_),
    .SUM(_00646_));
 sky130_fd_sc_hd__ha_1 _27711_ (.A(net393),
    .B(net387),
    .COUT(_13524_),
    .SUM(_00647_));
 sky130_fd_sc_hd__ha_1 _27712_ (.A(\count15_2[1] ),
    .B(net1133),
    .COUT(_13525_),
    .SUM(_00648_));
 sky130_fd_sc_hd__ha_1 _27713_ (.A(net471),
    .B(net466),
    .COUT(_13526_),
    .SUM(_00649_));
 sky130_fd_sc_hd__ha_4 _27714_ (.A(_00650_),
    .B(_13527_),
    .COUT(_13528_),
    .SUM(_00651_));
 sky130_fd_sc_hd__ha_4 _27715_ (.A(_00650_),
    .B(\count_1[2] ),
    .COUT(_13529_),
    .SUM(_13530_));
 sky130_fd_sc_hd__ha_4 _27716_ (.A(\count_1[1] ),
    .B(_13527_),
    .COUT(_13531_),
    .SUM(_13532_));
 sky130_fd_sc_hd__ha_4 _27717_ (.A(\count_1[1] ),
    .B(\count_1[2] ),
    .COUT(_13533_),
    .SUM(_13534_));
 sky130_fd_sc_hd__ha_4 _27718_ (.A(_00652_),
    .B(_13535_),
    .COUT(_13536_),
    .SUM(_00653_));
 sky130_fd_sc_hd__ha_4 _27719_ (.A(_00652_),
    .B(\count_2[2] ),
    .COUT(_13537_),
    .SUM(_13538_));
 sky130_fd_sc_hd__ha_4 _27720_ (.A(\count_2[1] ),
    .B(_13535_),
    .COUT(_13539_),
    .SUM(_13540_));
 sky130_fd_sc_hd__ha_4 _27721_ (.A(\count_2[1] ),
    .B(\count_2[2] ),
    .COUT(_13541_),
    .SUM(_13542_));
 sky130_fd_sc_hd__ha_2 _27722_ (.A(_00658_),
    .B(_13543_),
    .COUT(_13544_),
    .SUM(_13545_));
 sky130_fd_sc_hd__ha_1 _27723_ (.A(net1093),
    .B(\count2_1[2] ),
    .COUT(_13546_),
    .SUM(_00642_));
 sky130_fd_sc_hd__ha_1 _27724_ (.A(_13547_),
    .B(_13548_),
    .COUT(_13549_),
    .SUM(_13550_));
 sky130_fd_sc_hd__ha_1 _27725_ (.A(_13551_),
    .B(_13552_),
    .COUT(_13553_),
    .SUM(_13554_));
 sky130_fd_sc_hd__ha_4 _27726_ (.A(_13555_),
    .B(_13556_),
    .COUT(_13557_),
    .SUM(_13558_));
 sky130_fd_sc_hd__ha_1 _27727_ (.A(_13559_),
    .B(_13560_),
    .COUT(_13561_),
    .SUM(_13562_));
 sky130_fd_sc_hd__ha_1 _27728_ (.A(_13563_),
    .B(_13564_),
    .COUT(_13565_),
    .SUM(_13566_));
 sky130_fd_sc_hd__ha_2 _27729_ (.A(_13567_),
    .B(_13568_),
    .COUT(_13569_),
    .SUM(_13570_));
 sky130_fd_sc_hd__ha_1 _27730_ (.A(_13571_),
    .B(_13572_),
    .COUT(_13573_),
    .SUM(_13574_));
 sky130_fd_sc_hd__ha_4 _27731_ (.A(_13575_),
    .B(_13576_),
    .COUT(_13577_),
    .SUM(_13578_));
 sky130_fd_sc_hd__ha_4 _27732_ (.A(_13579_),
    .B(_13580_),
    .COUT(_13581_),
    .SUM(_13582_));
 sky130_fd_sc_hd__ha_4 _27733_ (.A(_13583_),
    .B(_13584_),
    .COUT(_13585_),
    .SUM(_13586_));
 sky130_fd_sc_hd__ha_1 _27734_ (.A(_13587_),
    .B(_13588_),
    .COUT(_13589_),
    .SUM(_13590_));
 sky130_fd_sc_hd__ha_1 _27735_ (.A(_13591_),
    .B(_13592_),
    .COUT(_13593_),
    .SUM(_13594_));
 sky130_fd_sc_hd__ha_4 _27736_ (.A(_13595_),
    .B(_13596_),
    .COUT(_13597_),
    .SUM(_13598_));
 sky130_fd_sc_hd__ha_1 _27737_ (.A(_13599_),
    .B(_13600_),
    .COUT(_13601_),
    .SUM(_13602_));
 sky130_fd_sc_hd__ha_2 _27738_ (.A(_13603_),
    .B(_13604_),
    .COUT(_13605_),
    .SUM(_13606_));
 sky130_fd_sc_hd__ha_4 _27739_ (.A(_13607_),
    .B(_13608_),
    .COUT(_13609_),
    .SUM(_13610_));
 sky130_fd_sc_hd__ha_1 _27740_ (.A(_13611_),
    .B(_13612_),
    .COUT(_13613_),
    .SUM(_13614_));
 sky130_fd_sc_hd__ha_4 _27741_ (.A(_13615_),
    .B(_13616_),
    .COUT(_13617_),
    .SUM(_13618_));
 sky130_fd_sc_hd__ha_4 _27742_ (.A(_13619_),
    .B(_13620_),
    .COUT(_13621_),
    .SUM(_13622_));
 sky130_fd_sc_hd__ha_4 _27743_ (.A(_13623_),
    .B(_13624_),
    .COUT(_13625_),
    .SUM(_13626_));
 sky130_fd_sc_hd__ha_4 _27744_ (.A(_13627_),
    .B(_13628_),
    .COUT(_13629_),
    .SUM(_13630_));
 sky130_fd_sc_hd__ha_1 _27745_ (.A(_13631_),
    .B(_13632_),
    .COUT(_13633_),
    .SUM(_13634_));
 sky130_fd_sc_hd__ha_1 _27746_ (.A(_13635_),
    .B(_13636_),
    .COUT(_13637_),
    .SUM(_13638_));
 sky130_fd_sc_hd__ha_4 _27747_ (.A(_13639_),
    .B(_13640_),
    .COUT(_13641_),
    .SUM(_13642_));
 sky130_fd_sc_hd__ha_2 _27748_ (.A(_13643_),
    .B(_13644_),
    .COUT(_13645_),
    .SUM(_13646_));
 sky130_fd_sc_hd__ha_2 _27749_ (.A(_13647_),
    .B(_13648_),
    .COUT(_13649_),
    .SUM(_13650_));
 sky130_fd_sc_hd__ha_1 _27750_ (.A(_13651_),
    .B(_13652_),
    .COUT(_13653_),
    .SUM(_13654_));
 sky130_fd_sc_hd__ha_1 _27751_ (.A(_13655_),
    .B(_13656_),
    .COUT(_13657_),
    .SUM(_13658_));
 sky130_fd_sc_hd__ha_1 _27752_ (.A(_13659_),
    .B(_13660_),
    .COUT(_13661_),
    .SUM(_13662_));
 sky130_fd_sc_hd__ha_1 _27753_ (.A(_13663_),
    .B(_13664_),
    .COUT(_13665_),
    .SUM(_13666_));
 sky130_fd_sc_hd__ha_2 _27754_ (.A(_13667_),
    .B(_13668_),
    .COUT(_12378_),
    .SUM(\hash.CA1.p4[1] ));
 sky130_fd_sc_hd__ha_1 _27755_ (.A(_12899_),
    .B(\hash.CA1.p4[1] ),
    .COUT(_13669_),
    .SUM(_13670_));
 sky130_fd_sc_hd__ha_1 _27756_ (.A(_12379_),
    .B(_12377_),
    .COUT(_13671_),
    .SUM(_13672_));
 sky130_fd_sc_hd__ha_1 _27757_ (.A(\hash.CA1.p4[2] ),
    .B(_13673_),
    .COUT(_13674_),
    .SUM(_13675_));
 sky130_fd_sc_hd__ha_1 _27758_ (.A(_12376_),
    .B(_13676_),
    .COUT(_13677_),
    .SUM(_13678_));
 sky130_fd_sc_hd__ha_1 _27759_ (.A(\hash.CA1.p4[3] ),
    .B(_13679_),
    .COUT(_13680_),
    .SUM(_13681_));
 sky130_fd_sc_hd__ha_1 _27760_ (.A(_13682_),
    .B(_12388_),
    .COUT(_13683_),
    .SUM(_13684_));
 sky130_fd_sc_hd__ha_4 _27761_ (.A(\hash.CA1.p4[4] ),
    .B(_13685_),
    .COUT(_13686_),
    .SUM(_13687_));
 sky130_fd_sc_hd__ha_1 _27762_ (.A(_12387_),
    .B(_13688_),
    .COUT(_13689_),
    .SUM(_13690_));
 sky130_fd_sc_hd__ha_4 _27763_ (.A(\hash.CA1.p4[5] ),
    .B(_13691_),
    .COUT(_13692_),
    .SUM(_13693_));
 sky130_fd_sc_hd__ha_1 _27764_ (.A(_13694_),
    .B(_12396_),
    .COUT(_13695_),
    .SUM(_13696_));
 sky130_fd_sc_hd__ha_4 _27765_ (.A(\hash.CA1.p4[6] ),
    .B(_13697_),
    .COUT(_13698_),
    .SUM(_13699_));
 sky130_fd_sc_hd__ha_1 _27766_ (.A(_12395_),
    .B(_13700_),
    .COUT(_13701_),
    .SUM(_13702_));
 sky130_fd_sc_hd__ha_1 _27767_ (.A(\hash.CA1.p4[7] ),
    .B(_13703_),
    .COUT(_13704_),
    .SUM(_13705_));
 sky130_fd_sc_hd__ha_1 _27768_ (.A(_13706_),
    .B(_13707_),
    .COUT(_13708_),
    .SUM(_13709_));
 sky130_fd_sc_hd__ha_1 _27769_ (.A(\hash.CA1.p4[8] ),
    .B(_13710_),
    .COUT(_13711_),
    .SUM(_13712_));
 sky130_fd_sc_hd__ha_2 _27770_ (.A(_13713_),
    .B(_12409_),
    .COUT(_13714_),
    .SUM(_13715_));
 sky130_fd_sc_hd__ha_1 _27771_ (.A(\hash.CA1.p4[9] ),
    .B(_13716_),
    .COUT(_13717_),
    .SUM(_13718_));
 sky130_fd_sc_hd__ha_4 _27772_ (.A(_12408_),
    .B(_12412_),
    .COUT(_13719_),
    .SUM(_13720_));
 sky130_fd_sc_hd__ha_1 _27773_ (.A(\hash.CA1.p4[10] ),
    .B(_13721_),
    .COUT(_13722_),
    .SUM(_13723_));
 sky130_fd_sc_hd__ha_4 _27774_ (.A(_12411_),
    .B(_13724_),
    .COUT(_13725_),
    .SUM(_13726_));
 sky130_fd_sc_hd__ha_2 _27775_ (.A(\hash.CA1.p4[11] ),
    .B(_13727_),
    .COUT(_13728_),
    .SUM(_13729_));
 sky130_fd_sc_hd__ha_4 _27776_ (.A(_13730_),
    .B(_13731_),
    .COUT(_13732_),
    .SUM(_13733_));
 sky130_fd_sc_hd__ha_4 _27777_ (.A(\hash.CA1.p4[12] ),
    .B(_13734_),
    .COUT(_13735_),
    .SUM(_13736_));
 sky130_fd_sc_hd__ha_1 _27778_ (.A(_13737_),
    .B(_12425_),
    .COUT(_13738_),
    .SUM(_13739_));
 sky130_fd_sc_hd__ha_4 _27779_ (.A(\hash.CA1.p4[13] ),
    .B(_13740_),
    .COUT(_13741_),
    .SUM(_13742_));
 sky130_fd_sc_hd__ha_1 _27780_ (.A(_12424_),
    .B(_13743_),
    .COUT(_13744_),
    .SUM(_13745_));
 sky130_fd_sc_hd__ha_2 _27781_ (.A(\hash.CA1.p4[14] ),
    .B(_13746_),
    .COUT(_13747_),
    .SUM(_13748_));
 sky130_fd_sc_hd__ha_1 _27782_ (.A(_13749_),
    .B(_13750_),
    .COUT(_13751_),
    .SUM(_13752_));
 sky130_fd_sc_hd__ha_2 _27783_ (.A(\hash.CA1.p4[15] ),
    .B(_13753_),
    .COUT(_13754_),
    .SUM(_13755_));
 sky130_fd_sc_hd__ha_1 _27784_ (.A(_13756_),
    .B(_13757_),
    .COUT(_13758_),
    .SUM(_13759_));
 sky130_fd_sc_hd__ha_2 _27785_ (.A(\hash.CA1.p4[16] ),
    .B(_13760_),
    .COUT(_13761_),
    .SUM(_13762_));
 sky130_fd_sc_hd__ha_1 _27786_ (.A(_13763_),
    .B(_13764_),
    .COUT(_13765_),
    .SUM(_13766_));
 sky130_fd_sc_hd__ha_1 _27787_ (.A(\hash.CA1.p4[17] ),
    .B(_13767_),
    .COUT(_13768_),
    .SUM(_13769_));
 sky130_fd_sc_hd__ha_1 _27788_ (.A(_13770_),
    .B(_12448_),
    .COUT(_13771_),
    .SUM(_13772_));
 sky130_fd_sc_hd__ha_1 _27789_ (.A(\hash.CA1.p4[18] ),
    .B(_13773_),
    .COUT(_13774_),
    .SUM(_13775_));
 sky130_fd_sc_hd__ha_1 _27790_ (.A(_12447_),
    .B(_12451_),
    .COUT(_13776_),
    .SUM(_13777_));
 sky130_fd_sc_hd__ha_1 _27791_ (.A(\hash.CA1.p4[19] ),
    .B(_13778_),
    .COUT(_13779_),
    .SUM(_13780_));
 sky130_fd_sc_hd__ha_4 _27792_ (.A(_12450_),
    .B(_12454_),
    .COUT(_13781_),
    .SUM(_13782_));
 sky130_fd_sc_hd__ha_1 _27793_ (.A(\hash.CA1.p4[20] ),
    .B(_13783_),
    .COUT(_13784_),
    .SUM(_13785_));
 sky130_fd_sc_hd__ha_4 _27794_ (.A(_12453_),
    .B(_12457_),
    .COUT(_13786_),
    .SUM(_13787_));
 sky130_fd_sc_hd__ha_4 _27795_ (.A(\hash.CA1.p4[21] ),
    .B(_13788_),
    .COUT(_13789_),
    .SUM(_13790_));
 sky130_fd_sc_hd__ha_1 _27796_ (.A(_12456_),
    .B(_12460_),
    .COUT(_13791_),
    .SUM(_13792_));
 sky130_fd_sc_hd__ha_1 _27797_ (.A(\hash.CA1.p4[22] ),
    .B(_13793_),
    .COUT(_13794_),
    .SUM(_13795_));
 sky130_fd_sc_hd__ha_1 _27798_ (.A(_12459_),
    .B(_13796_),
    .COUT(_13797_),
    .SUM(_13798_));
 sky130_fd_sc_hd__ha_1 _27799_ (.A(\hash.CA1.p4[23] ),
    .B(_13799_),
    .COUT(_13800_),
    .SUM(_13801_));
 sky130_fd_sc_hd__ha_1 _27800_ (.A(_13802_),
    .B(_13803_),
    .COUT(_13804_),
    .SUM(_13805_));
 sky130_fd_sc_hd__ha_1 _27801_ (.A(\hash.CA1.p4[24] ),
    .B(_13806_),
    .COUT(_13807_),
    .SUM(_13808_));
 sky130_fd_sc_hd__ha_1 _27802_ (.A(_13809_),
    .B(_13810_),
    .COUT(_13811_),
    .SUM(_13812_));
 sky130_fd_sc_hd__ha_1 _27803_ (.A(\hash.CA1.p4[25] ),
    .B(_13813_),
    .COUT(_13814_),
    .SUM(_13815_));
 sky130_fd_sc_hd__ha_1 _27804_ (.A(_13816_),
    .B(_13817_),
    .COUT(_13818_),
    .SUM(_13819_));
 sky130_fd_sc_hd__ha_4 _27805_ (.A(\hash.CA1.p4[26] ),
    .B(_06287_),
    .COUT(_13821_),
    .SUM(_13822_));
 sky130_fd_sc_hd__ha_2 _27806_ (.A(_13823_),
    .B(_13824_),
    .COUT(_13825_),
    .SUM(_13826_));
 sky130_fd_sc_hd__ha_4 _27807_ (.A(\hash.CA1.p4[27] ),
    .B(_13827_),
    .COUT(_13828_),
    .SUM(_13829_));
 sky130_fd_sc_hd__ha_1 _27808_ (.A(_13830_),
    .B(_13831_),
    .COUT(_13832_),
    .SUM(_13833_));
 sky130_fd_sc_hd__ha_1 _27809_ (.A(\hash.CA1.p4[28] ),
    .B(_13834_),
    .COUT(_13835_),
    .SUM(_13836_));
 sky130_fd_sc_hd__ha_4 _27810_ (.A(_13837_),
    .B(_12493_),
    .COUT(_13838_),
    .SUM(_13839_));
 sky130_fd_sc_hd__ha_1 _27811_ (.A(\hash.CA1.p4[29] ),
    .B(_13840_),
    .COUT(_13841_),
    .SUM(_13842_));
 sky130_fd_sc_hd__ha_1 _27812_ (.A(_12492_),
    .B(_12496_),
    .COUT(_13843_),
    .SUM(_13844_));
 sky130_fd_sc_hd__ha_1 _27813_ (.A(\hash.CA1.p4[30] ),
    .B(_13845_),
    .COUT(_13846_),
    .SUM(_13847_));
 sky130_fd_sc_hd__ha_1 _27814_ (.A(_12653_),
    .B(_12505_),
    .COUT(_13848_),
    .SUM(_11578_));
 sky130_fd_sc_hd__ha_4 _27815_ (.A(_00843_),
    .B(_12368_),
    .COUT(_13849_),
    .SUM(_13850_));
 sky130_fd_sc_hd__ha_4 _27816_ (.A(_00813_),
    .B(_13851_),
    .COUT(_13852_),
    .SUM(_13853_));
 sky130_fd_sc_hd__ha_4 _27817_ (.A(_13854_),
    .B(_00781_),
    .COUT(_13855_),
    .SUM(_13856_));
 sky130_fd_sc_hd__ha_1 _27818_ (.A(_12657_),
    .B(_13857_),
    .COUT(_13858_),
    .SUM(_11577_));
 sky130_fd_sc_hd__ha_4 _27819_ (.A(_12899_),
    .B(_13673_),
    .COUT(_13859_),
    .SUM(_11576_));
 sky130_fd_sc_hd__ha_4 _27820_ (.A(\hash.CA1.b[1] ),
    .B(\hash.CA1.b[0] ),
    .COUT(_13860_),
    .SUM(_11575_));
 sky130_fd_sc_hd__ha_4 _27821_ (.A(\hash.CA1.k_i1[0] ),
    .B(\hash.CA1.w_i1[0] ),
    .COUT(_12497_),
    .SUM(_12654_));
 sky130_fd_sc_hd__ha_4 _27822_ (.A(_13862_),
    .B(_13861_),
    .COUT(_12500_),
    .SUM(_12887_));
 sky130_fd_sc_hd__ha_1 _27823_ (.A(\hash.CA1.k_i1[1] ),
    .B(\hash.CA1.w_i1[1] ),
    .COUT(_13863_),
    .SUM(_13864_));
 sky130_fd_sc_hd__ha_1 _27824_ (.A(_12501_),
    .B(_12502_),
    .COUT(_13865_),
    .SUM(_13866_));
 sky130_fd_sc_hd__ha_1 _27825_ (.A(\hash.CA1.k_i1[2] ),
    .B(\hash.CA1.w_i1[2] ),
    .COUT(_13867_),
    .SUM(_13868_));
 sky130_fd_sc_hd__ha_1 _27826_ (.A(_13869_),
    .B(_13870_),
    .COUT(_13871_),
    .SUM(_13872_));
 sky130_fd_sc_hd__ha_1 _27827_ (.A(_12506_),
    .B(_12512_),
    .COUT(_13873_),
    .SUM(_13874_));
 sky130_fd_sc_hd__ha_1 _27828_ (.A(\hash.CA1.k_i1[3] ),
    .B(\hash.CA1.w_i1[3] ),
    .COUT(_13875_),
    .SUM(_13876_));
 sky130_fd_sc_hd__ha_4 _27829_ (.A(_13877_),
    .B(_13878_),
    .COUT(_13879_),
    .SUM(_13880_));
 sky130_fd_sc_hd__ha_4 _27830_ (.A(_12511_),
    .B(_13881_),
    .COUT(_13882_),
    .SUM(_13883_));
 sky130_fd_sc_hd__ha_1 _27831_ (.A(\hash.CA1.k_i1[4] ),
    .B(\hash.CA1.w_i1[4] ),
    .COUT(_13884_),
    .SUM(_13885_));
 sky130_fd_sc_hd__ha_4 _27832_ (.A(_13887_),
    .B(_13886_),
    .COUT(_13888_),
    .SUM(_13889_));
 sky130_fd_sc_hd__ha_1 _27833_ (.A(_13890_),
    .B(_13891_),
    .COUT(_13892_),
    .SUM(_13893_));
 sky130_fd_sc_hd__ha_4 _27834_ (.A(\hash.CA1.k_i1[5] ),
    .B(\hash.CA1.w_i1[5] ),
    .COUT(_13894_),
    .SUM(_13895_));
 sky130_fd_sc_hd__ha_2 _27835_ (.A(_13896_),
    .B(_13897_),
    .COUT(_13898_),
    .SUM(_13899_));
 sky130_fd_sc_hd__ha_1 _27836_ (.A(_13900_),
    .B(_12527_),
    .COUT(_13901_),
    .SUM(_13902_));
 sky130_fd_sc_hd__ha_1 _27837_ (.A(\hash.CA1.k_i1[6] ),
    .B(\hash.CA1.w_i1[6] ),
    .COUT(_13903_),
    .SUM(_13904_));
 sky130_fd_sc_hd__ha_2 _27838_ (.A(_13905_),
    .B(_13906_),
    .COUT(_13907_),
    .SUM(_13908_));
 sky130_fd_sc_hd__ha_4 _27839_ (.A(_12526_),
    .B(_12532_),
    .COUT(_13909_),
    .SUM(_13910_));
 sky130_fd_sc_hd__ha_2 _27840_ (.A(\hash.CA1.k_i1[7] ),
    .B(\hash.CA1.w_i1[7] ),
    .COUT(_13911_),
    .SUM(_13912_));
 sky130_fd_sc_hd__ha_4 _27841_ (.A(_13913_),
    .B(_13914_),
    .COUT(_13915_),
    .SUM(_13916_));
 sky130_fd_sc_hd__ha_4 _27842_ (.A(_12531_),
    .B(_12537_),
    .COUT(_13917_),
    .SUM(_13918_));
 sky130_fd_sc_hd__ha_1 _27843_ (.A(\hash.CA1.k_i1[8] ),
    .B(\hash.CA1.w_i1[8] ),
    .COUT(_13919_),
    .SUM(_13920_));
 sky130_fd_sc_hd__ha_4 _27844_ (.A(_13921_),
    .B(_13922_),
    .COUT(_13923_),
    .SUM(_13924_));
 sky130_fd_sc_hd__ha_4 _27845_ (.A(_12536_),
    .B(_13925_),
    .COUT(_13926_),
    .SUM(_13927_));
 sky130_fd_sc_hd__ha_1 _27846_ (.A(\hash.CA1.k_i1[9] ),
    .B(\hash.CA1.w_i1[9] ),
    .COUT(_13928_),
    .SUM(_13929_));
 sky130_fd_sc_hd__ha_1 _27847_ (.A(_13930_),
    .B(_13931_),
    .COUT(_13932_),
    .SUM(_13933_));
 sky130_fd_sc_hd__ha_4 _27848_ (.A(_12547_),
    .B(_13934_),
    .COUT(_13935_),
    .SUM(_13936_));
 sky130_fd_sc_hd__ha_1 _27849_ (.A(\hash.CA1.k_i1[10] ),
    .B(\hash.CA1.w_i1[10] ),
    .COUT(_13937_),
    .SUM(_13938_));
 sky130_fd_sc_hd__ha_1 _27850_ (.A(_13939_),
    .B(_13940_),
    .COUT(_13941_),
    .SUM(_13942_));
 sky130_fd_sc_hd__ha_4 _27851_ (.A(_13943_),
    .B(_12546_),
    .COUT(_13944_),
    .SUM(_13945_));
 sky130_fd_sc_hd__ha_1 _27852_ (.A(\hash.CA1.k_i1[11] ),
    .B(\hash.CA1.w_i1[11] ),
    .COUT(_13946_),
    .SUM(_13947_));
 sky130_fd_sc_hd__ha_4 _27853_ (.A(_13948_),
    .B(_13949_),
    .COUT(_13950_),
    .SUM(_13951_));
 sky130_fd_sc_hd__ha_4 _27854_ (.A(_13952_),
    .B(_13953_),
    .COUT(_13954_),
    .SUM(_13955_));
 sky130_fd_sc_hd__ha_1 _27855_ (.A(\hash.CA1.k_i1[12] ),
    .B(\hash.CA1.w_i1[12] ),
    .COUT(_13956_),
    .SUM(_13957_));
 sky130_fd_sc_hd__ha_1 _27856_ (.A(_13958_),
    .B(_13959_),
    .COUT(_13960_),
    .SUM(_13961_));
 sky130_fd_sc_hd__ha_4 _27857_ (.A(_13962_),
    .B(_12562_),
    .COUT(_13963_),
    .SUM(_13964_));
 sky130_fd_sc_hd__ha_1 _27858_ (.A(\hash.CA1.k_i1[13] ),
    .B(\hash.CA1.w_i1[13] ),
    .COUT(_13965_),
    .SUM(_13966_));
 sky130_fd_sc_hd__ha_4 _27859_ (.A(_13967_),
    .B(_13968_),
    .COUT(_13969_),
    .SUM(_13970_));
 sky130_fd_sc_hd__ha_2 _27860_ (.A(_12561_),
    .B(_12567_),
    .COUT(_13971_),
    .SUM(_13972_));
 sky130_fd_sc_hd__ha_4 _27861_ (.A(\hash.CA1.k_i1[14] ),
    .B(\hash.CA1.w_i1[14] ),
    .COUT(_13973_),
    .SUM(_13974_));
 sky130_fd_sc_hd__ha_4 _27862_ (.A(_13975_),
    .B(_13976_),
    .COUT(_13977_),
    .SUM(_13978_));
 sky130_fd_sc_hd__ha_4 _27863_ (.A(_13979_),
    .B(_12566_),
    .COUT(_13980_),
    .SUM(_13981_));
 sky130_fd_sc_hd__ha_1 _27864_ (.A(\hash.CA1.k_i1[15] ),
    .B(\hash.CA1.w_i1[15] ),
    .COUT(_13982_),
    .SUM(_13983_));
 sky130_fd_sc_hd__ha_4 _27865_ (.A(_13984_),
    .B(_13985_),
    .COUT(_13986_),
    .SUM(_13987_));
 sky130_fd_sc_hd__ha_4 _27866_ (.A(_13988_),
    .B(_13989_),
    .COUT(_13990_),
    .SUM(_13991_));
 sky130_fd_sc_hd__ha_1 _27867_ (.A(\hash.CA1.k_i1[16] ),
    .B(\hash.CA1.w_i1[16] ),
    .COUT(_13992_),
    .SUM(_13993_));
 sky130_fd_sc_hd__ha_4 _27868_ (.A(_13994_),
    .B(_13995_),
    .COUT(_13996_),
    .SUM(_13997_));
 sky130_fd_sc_hd__ha_4 _27869_ (.A(_13998_),
    .B(_12582_),
    .COUT(_13999_),
    .SUM(_14000_));
 sky130_fd_sc_hd__ha_1 _27870_ (.A(\hash.CA1.k_i1[17] ),
    .B(\hash.CA1.w_i1[17] ),
    .COUT(_14001_),
    .SUM(_14002_));
 sky130_fd_sc_hd__ha_4 _27871_ (.A(_14003_),
    .B(_14004_),
    .COUT(_14005_),
    .SUM(_14006_));
 sky130_fd_sc_hd__ha_4 _27872_ (.A(_12581_),
    .B(_12587_),
    .COUT(_14007_),
    .SUM(_14008_));
 sky130_fd_sc_hd__ha_1 _27873_ (.A(\hash.CA1.k_i1[18] ),
    .B(\hash.CA1.w_i1[18] ),
    .COUT(_14009_),
    .SUM(_14010_));
 sky130_fd_sc_hd__ha_2 _27874_ (.A(_14011_),
    .B(_14012_),
    .COUT(_14013_),
    .SUM(_14014_));
 sky130_fd_sc_hd__ha_4 _27875_ (.A(_12586_),
    .B(_12592_),
    .COUT(_14015_),
    .SUM(_14016_));
 sky130_fd_sc_hd__ha_1 _27876_ (.A(\hash.CA1.k_i1[19] ),
    .B(\hash.CA1.w_i1[19] ),
    .COUT(_14017_),
    .SUM(_14018_));
 sky130_fd_sc_hd__ha_1 _27877_ (.A(_14019_),
    .B(_14020_),
    .COUT(_14021_),
    .SUM(_14022_));
 sky130_fd_sc_hd__ha_4 _27878_ (.A(_12591_),
    .B(_12597_),
    .COUT(_14023_),
    .SUM(_14024_));
 sky130_fd_sc_hd__ha_1 _27879_ (.A(\hash.CA1.k_i1[20] ),
    .B(\hash.CA1.w_i1[20] ),
    .COUT(_14025_),
    .SUM(_14026_));
 sky130_fd_sc_hd__ha_1 _27880_ (.A(_14027_),
    .B(_14028_),
    .COUT(_14029_),
    .SUM(_14030_));
 sky130_fd_sc_hd__ha_2 _27881_ (.A(_12596_),
    .B(_12602_),
    .COUT(_14031_),
    .SUM(_14032_));
 sky130_fd_sc_hd__ha_2 _27882_ (.A(\hash.CA1.k_i1[21] ),
    .B(\hash.CA1.w_i1[21] ),
    .COUT(_14033_),
    .SUM(_14034_));
 sky130_fd_sc_hd__ha_1 _27883_ (.A(_14035_),
    .B(_14036_),
    .COUT(_14037_),
    .SUM(_14038_));
 sky130_fd_sc_hd__ha_1 _27884_ (.A(_12601_),
    .B(_14039_),
    .COUT(_14040_),
    .SUM(_14041_));
 sky130_fd_sc_hd__ha_4 _27885_ (.A(\hash.CA1.k_i1[22] ),
    .B(\hash.CA1.w_i1[22] ),
    .COUT(_14042_),
    .SUM(_14043_));
 sky130_fd_sc_hd__ha_1 _27886_ (.A(_14044_),
    .B(_14045_),
    .COUT(_14046_),
    .SUM(_14047_));
 sky130_fd_sc_hd__ha_1 _27887_ (.A(_14048_),
    .B(_14049_),
    .COUT(_14050_),
    .SUM(_14051_));
 sky130_fd_sc_hd__ha_1 _27888_ (.A(\hash.CA1.k_i1[23] ),
    .B(\hash.CA1.w_i1[23] ),
    .COUT(_14052_),
    .SUM(_14053_));
 sky130_fd_sc_hd__ha_2 _27889_ (.A(_14054_),
    .B(_14055_),
    .COUT(_14056_),
    .SUM(_14057_));
 sky130_fd_sc_hd__ha_4 _27890_ (.A(_14058_),
    .B(_14059_),
    .COUT(_14060_),
    .SUM(_14061_));
 sky130_fd_sc_hd__ha_1 _27891_ (.A(\hash.CA1.k_i1[24] ),
    .B(\hash.CA1.w_i1[24] ),
    .COUT(_14062_),
    .SUM(_14063_));
 sky130_fd_sc_hd__ha_4 _27892_ (.A(_14064_),
    .B(_14065_),
    .COUT(_14066_),
    .SUM(_14067_));
 sky130_fd_sc_hd__ha_4 _27893_ (.A(_14068_),
    .B(_14069_),
    .COUT(_14070_),
    .SUM(_14071_));
 sky130_fd_sc_hd__ha_2 _27894_ (.A(\hash.CA1.k_i1[25] ),
    .B(\hash.CA1.w_i1[25] ),
    .COUT(_14072_),
    .SUM(_14073_));
 sky130_fd_sc_hd__ha_1 _27895_ (.A(_14074_),
    .B(_14075_),
    .COUT(_14076_),
    .SUM(_14077_));
 sky130_fd_sc_hd__ha_4 _27896_ (.A(_14078_),
    .B(_14079_),
    .COUT(_14080_),
    .SUM(_14081_));
 sky130_fd_sc_hd__ha_2 _27897_ (.A(\hash.CA1.k_i1[26] ),
    .B(\hash.CA1.w_i1[26] ),
    .COUT(_14082_),
    .SUM(_14083_));
 sky130_fd_sc_hd__ha_2 _27898_ (.A(_14084_),
    .B(_14085_),
    .COUT(_14086_),
    .SUM(_14087_));
 sky130_fd_sc_hd__ha_2 _27899_ (.A(_14088_),
    .B(_12632_),
    .COUT(_14089_),
    .SUM(_14090_));
 sky130_fd_sc_hd__ha_1 _27900_ (.A(\hash.CA1.k_i1[27] ),
    .B(\hash.CA1.w_i1[27] ),
    .COUT(_14091_),
    .SUM(_14092_));
 sky130_fd_sc_hd__ha_4 _27901_ (.A(_14093_),
    .B(_14094_),
    .COUT(_14095_),
    .SUM(_14096_));
 sky130_fd_sc_hd__ha_2 _27902_ (.A(_12631_),
    .B(_14097_),
    .COUT(_14098_),
    .SUM(_14099_));
 sky130_fd_sc_hd__ha_1 _27903_ (.A(\hash.CA1.k_i1[28] ),
    .B(\hash.CA1.w_i1[28] ),
    .COUT(_14100_),
    .SUM(_14101_));
 sky130_fd_sc_hd__ha_1 _27904_ (.A(_14102_),
    .B(_14103_),
    .COUT(_14104_),
    .SUM(_14105_));
 sky130_fd_sc_hd__ha_2 _27905_ (.A(_14106_),
    .B(_14107_),
    .COUT(_14108_),
    .SUM(_14109_));
 sky130_fd_sc_hd__ha_1 _27906_ (.A(\hash.CA1.k_i1[29] ),
    .B(\hash.CA1.w_i1[29] ),
    .COUT(_14110_),
    .SUM(_14111_));
 sky130_fd_sc_hd__ha_1 _27907_ (.A(_14112_),
    .B(_14113_),
    .COUT(_14114_),
    .SUM(_14115_));
 sky130_fd_sc_hd__ha_1 _27908_ (.A(_14116_),
    .B(_12647_),
    .COUT(_14117_),
    .SUM(_14118_));
 sky130_fd_sc_hd__ha_1 _27909_ (.A(\hash.CA1.k_i1[30] ),
    .B(\hash.CA1.w_i1[30] ),
    .COUT(_14119_),
    .SUM(_14120_));
 sky130_fd_sc_hd__ha_1 _27910_ (.A(_14121_),
    .B(_14122_),
    .COUT(_14123_),
    .SUM(_14124_));
 sky130_fd_sc_hd__ha_1 _27911_ (.A(_12646_),
    .B(_14125_),
    .COUT(_14126_),
    .SUM(_14127_));
 sky130_fd_sc_hd__ha_1 _27912_ (.A(_14128_),
    .B(_14129_),
    .COUT(_14130_),
    .SUM(_14131_));
 sky130_fd_sc_hd__ha_1 _27913_ (.A(_14132_),
    .B(_14133_),
    .COUT(_14134_),
    .SUM(_14135_));
 sky130_fd_sc_hd__ha_4 _27914_ (.A(_14136_),
    .B(_14137_),
    .COUT(_14138_),
    .SUM(_14139_));
 sky130_fd_sc_hd__ha_4 _27915_ (.A(_14140_),
    .B(_14141_),
    .COUT(_14142_),
    .SUM(_14143_));
 sky130_fd_sc_hd__ha_4 _27916_ (.A(_14144_),
    .B(_14145_),
    .COUT(_14146_),
    .SUM(_14147_));
 sky130_fd_sc_hd__ha_4 _27917_ (.A(_14148_),
    .B(_14149_),
    .COUT(_14150_),
    .SUM(_14151_));
 sky130_fd_sc_hd__ha_1 _27918_ (.A(_14152_),
    .B(_14153_),
    .COUT(_14154_),
    .SUM(_14155_));
 sky130_fd_sc_hd__ha_4 _27919_ (.A(_14156_),
    .B(_12722_),
    .COUT(_14157_),
    .SUM(_14158_));
 sky130_fd_sc_hd__ha_4 _27920_ (.A(_12730_),
    .B(_12721_),
    .COUT(_14159_),
    .SUM(_14160_));
 sky130_fd_sc_hd__ha_2 _27921_ (.A(_12729_),
    .B(_12739_),
    .COUT(_14161_),
    .SUM(_14162_));
 sky130_fd_sc_hd__ha_4 _27922_ (.A(_12738_),
    .B(_12745_),
    .COUT(_14163_),
    .SUM(_14164_));
 sky130_fd_sc_hd__ha_2 _27923_ (.A(_12744_),
    .B(_12751_),
    .COUT(_14165_),
    .SUM(_14166_));
 sky130_fd_sc_hd__ha_2 _27924_ (.A(_12750_),
    .B(_12758_),
    .COUT(_14167_),
    .SUM(_14168_));
 sky130_fd_sc_hd__ha_2 _27925_ (.A(_12757_),
    .B(_12766_),
    .COUT(_14169_),
    .SUM(_14170_));
 sky130_fd_sc_hd__ha_1 _27926_ (.A(_12765_),
    .B(_12773_),
    .COUT(_14171_),
    .SUM(_14172_));
 sky130_fd_sc_hd__ha_1 _27927_ (.A(_12772_),
    .B(_12779_),
    .COUT(_14173_),
    .SUM(_14174_));
 sky130_fd_sc_hd__ha_4 _27928_ (.A(_12778_),
    .B(_12785_),
    .COUT(_14175_),
    .SUM(_14176_));
 sky130_fd_sc_hd__ha_2 _27929_ (.A(_12784_),
    .B(_12791_),
    .COUT(_14177_),
    .SUM(_14178_));
 sky130_fd_sc_hd__ha_4 _27930_ (.A(_12790_),
    .B(_12800_),
    .COUT(_14179_),
    .SUM(_14180_));
 sky130_fd_sc_hd__ha_2 _27931_ (.A(_12799_),
    .B(_12809_),
    .COUT(_14181_),
    .SUM(_14182_));
 sky130_fd_sc_hd__ha_1 _27932_ (.A(_12808_),
    .B(_12816_),
    .COUT(_14183_),
    .SUM(_14184_));
 sky130_fd_sc_hd__ha_4 _27933_ (.A(_12815_),
    .B(_12825_),
    .COUT(_14185_),
    .SUM(_14186_));
 sky130_fd_sc_hd__ha_4 _27934_ (.A(_12824_),
    .B(_12832_),
    .COUT(_14187_),
    .SUM(_14188_));
 sky130_fd_sc_hd__ha_4 _27935_ (.A(_12831_),
    .B(_12841_),
    .COUT(_14189_),
    .SUM(_14190_));
 sky130_fd_sc_hd__ha_4 _27936_ (.A(_12840_),
    .B(_12847_),
    .COUT(_14191_),
    .SUM(_14192_));
 sky130_fd_sc_hd__ha_4 _27937_ (.A(_12846_),
    .B(_12855_),
    .COUT(_14193_),
    .SUM(_14194_));
 sky130_fd_sc_hd__ha_1 _27938_ (.A(_12854_),
    .B(_12863_),
    .COUT(_14195_),
    .SUM(_14196_));
 sky130_fd_sc_hd__ha_1 _27939_ (.A(_12862_),
    .B(_12869_),
    .COUT(_14197_),
    .SUM(_14198_));
 sky130_fd_sc_hd__ha_1 _27940_ (.A(_12868_),
    .B(_14199_),
    .COUT(_14200_),
    .SUM(_14201_));
 sky130_fd_sc_hd__ha_1 _27941_ (.A(_14202_),
    .B(_14203_),
    .COUT(_14204_),
    .SUM(\hash.CA1.p1[0] ));
 sky130_fd_sc_hd__ha_1 _27942_ (.A(_12656_),
    .B(_12887_),
    .COUT(_14205_),
    .SUM(\hash.CA1.p2[0] ));
 sky130_fd_sc_hd__ha_1 _27943_ (.A(_14205_),
    .B(_14206_),
    .COUT(_14207_),
    .SUM(\hash.CA1.p2[1] ));
 sky130_fd_sc_hd__ha_1 _27944_ (.A(_12888_),
    .B(_12507_),
    .COUT(_14208_),
    .SUM(\hash.CA1.p3[1] ));
 sky130_fd_sc_hd__ha_1 _27945_ (.A(\hash.CA1.c[0] ),
    .B(\hash.CA1.p4[0] ),
    .COUT(_12898_),
    .SUM(\hash.CA1.p5[0] ));
 sky130_fd_sc_hd__dfxtp_1 \count15_1[1]$_SDFF_PP0_  (.D(_00907_),
    .Q(\count15_1[1] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_4 \count15_1[2]$_SDFF_PP0_  (.D(_00908_),
    .Q(\count15_1[2] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 \count15_1[3]$_SDFF_PP0_  (.D(_00909_),
    .Q(\count15_1[3] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_1 \count15_1[4]$_SDFF_PP0_  (.D(_00910_),
    .Q(\count15_1[4] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_2 \count15_1[5]$_SDFF_PP0_  (.D(_00911_),
    .Q(\count15_1[5] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__dfxtp_2 \count15_2[1]$_SDFF_PP1_  (.D(_00912_),
    .Q(\count15_2[1] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_4 \count15_2[2]$_SDFF_PP0_  (.D(_00913_),
    .Q(\count15_2[2] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_2 \count15_2[3]$_SDFF_PP0_  (.D(_00914_),
    .Q(\count15_2[3] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \count15_2[4]$_SDFF_PP0_  (.D(_00915_),
    .Q(\count15_2[4] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 \count15_2[5]$_SDFF_PP0_  (.D(_00916_),
    .Q(\count15_2[5] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \count16_1[1]$_SDFF_PP0_  (.D(_00917_),
    .Q(\count16_1[1] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_2 \count16_1[2]$_SDFF_PP0_  (.D(_00918_),
    .Q(\count16_1[2] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \count16_1[3]$_SDFF_PP0_  (.D(_00919_),
    .Q(\count16_1[3] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \count16_1[4]$_SDFF_PP0_  (.D(_00920_),
    .Q(\count16_1[4] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 \count16_1[5]$_SDFF_PP0_  (.D(_00921_),
    .Q(\count16_1[5] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \count16_2[1]$_SDFF_PP0_  (.D(_00922_),
    .Q(\count16_2[1] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_2 \count16_2[2]$_SDFF_PP0_  (.D(_00923_),
    .Q(\count16_2[2] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_2 \count16_2[3]$_SDFF_PP0_  (.D(_00924_),
    .Q(\count16_2[3] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \count16_2[4]$_SDFF_PP0_  (.D(_00925_),
    .Q(\count16_2[4] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 \count16_2[5]$_SDFF_PP0_  (.D(_00926_),
    .Q(\count16_2[5] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_1[1]$_SDFF_PP1_  (.D(_00927_),
    .Q(\count2_1[1] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_4 \count2_1[2]$_SDFF_PP1_  (.D(_00928_),
    .Q(\count2_1[2] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_1[3]$_SDFF_PP1_  (.D(_00929_),
    .Q(\count2_1[3] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_1[4]$_SDFF_PP0_  (.D(_00930_),
    .Q(\count2_1[4] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_1[5]$_SDFF_PP0_  (.D(_00931_),
    .Q(\count2_1[5] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__dfxtp_4 \count2_2[1]$_SDFF_PP1_  (.D(_00932_),
    .Q(\count2_2[1] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_2[2]$_SDFF_PP1_  (.D(_00933_),
    .Q(\count2_2[2] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_2[3]$_SDFF_PP1_  (.D(_00934_),
    .Q(\count2_2[3] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_2[4]$_SDFF_PP0_  (.D(_00935_),
    .Q(\count2_2[4] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__dfxtp_1 \count2_2[5]$_SDFF_PP0_  (.D(_00936_),
    .Q(\count2_2[5] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_2 \count7_1[1]$_SDFF_PP0_  (.D(_00937_),
    .Q(\count7_1[1] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_1[2]$_SDFF_PP0_  (.D(_00938_),
    .Q(\count7_1[2] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_1[3]$_SDFF_PP1_  (.D(_00939_),
    .Q(\count7_1[3] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_1[4]$_SDFF_PP0_  (.D(_00940_),
    .Q(\count7_1[4] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__dfxtp_2 \count7_1[5]$_SDFF_PP0_  (.D(_00941_),
    .Q(\count7_1[5] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_2[1]$_SDFF_PP1_  (.D(_00942_),
    .Q(\count7_2[1] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_2[2]$_SDFF_PP0_  (.D(_00943_),
    .Q(\count7_2[2] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_2[3]$_SDFF_PP1_  (.D(_00944_),
    .Q(\count7_2[3] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_2[4]$_SDFF_PP0_  (.D(_00945_),
    .Q(\count7_2[4] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__dfxtp_1 \count7_2[5]$_SDFF_PP0_  (.D(_00946_),
    .Q(\count7_2[5] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_1[1]$_SDFFE_PP0N_  (.D(_00947_),
    .Q(\count_1[1] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_1[2]$_SDFFE_PP0N_  (.D(_00948_),
    .Q(\count_1[2] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_1[3]$_SDFFE_PP0N_  (.D(_00949_),
    .Q(\count_1[3] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_1[4]$_SDFFE_PP1N_  (.D(_00950_),
    .Q(\count_1[4] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_1[5]$_SDFFE_PP0N_  (.D(_00951_),
    .Q(\count_1[5] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[1]$_SDFFE_PP0N_  (.D(_00952_),
    .Q(\count_2[1] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[2]$_SDFFE_PP0N_  (.D(_00953_),
    .Q(\count_2[2] ),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[3]$_SDFFE_PP0N_  (.D(_00954_),
    .Q(\count_2[3] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[4]$_SDFFE_PP1N_  (.D(_00955_),
    .Q(\count_2[4] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[5]$_SDFFE_PP0N_  (.D(_00956_),
    .Q(\count_2[5] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_2[6]$_SDFFE_PP0N_  (.D(_00957_),
    .Q(\count_2[6] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash1[1]$_SDFFE_PP0N_  (.D(_00958_),
    .Q(\count_hash1[1] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash1[2]$_SDFFE_PP0N_  (.D(_00959_),
    .Q(\count_hash1[2] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash1[3]$_SDFFE_PP0N_  (.D(_00960_),
    .Q(\count_hash1[3] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash1[4]$_SDFFE_PP0N_  (.D(_00961_),
    .Q(\count_hash1[4] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash1[5]$_SDFFE_PP0N_  (.D(_00962_),
    .Q(\count_hash1[5] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash1[6]$_SDFFE_PP0N_  (.D(_00963_),
    .Q(\count_hash1[6] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash2[1]$_SDFFE_PP0N_  (.D(_00964_),
    .Q(\count_hash2[1] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash2[2]$_SDFFE_PP0N_  (.D(_00965_),
    .Q(\count_hash2[2] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash2[3]$_SDFFE_PP0N_  (.D(_00966_),
    .Q(\count_hash2[3] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash2[4]$_SDFFE_PP0N_  (.D(_00967_),
    .Q(\count_hash2[4] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 \count_hash2[5]$_SDFFE_PP0N_  (.D(_00968_),
    .Q(\count_hash2[5] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__edfxtp_1 \done$_DFFE_PN_  (.D(_00128_),
    .DE(_09731_),
    .Q(done),
    .CLK(clknet_leaf_55_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[0]$_DFF_P_  (.D(\hash.CA1.S0.X[0] ),
    .Q(\hash.CA2.a_dash[0] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[10]$_DFF_P_  (.D(\hash.CA1.S0.X[10] ),
    .Q(\hash.CA2.a_dash[10] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[11]$_DFF_P_  (.D(\hash.CA1.S0.X[11] ),
    .Q(\hash.CA2.a_dash[11] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[12]$_DFF_P_  (.D(\hash.CA1.S0.X[12] ),
    .Q(\hash.CA2.a_dash[12] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[13]$_DFF_P_  (.D(\hash.CA1.S0.X[13] ),
    .Q(\hash.CA2.a_dash[13] ),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[14]$_DFF_P_  (.D(\hash.CA1.S0.X[14] ),
    .Q(\hash.CA2.a_dash[14] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[15]$_DFF_P_  (.D(\hash.CA1.S0.X[15] ),
    .Q(\hash.CA2.a_dash[15] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[16]$_DFF_P_  (.D(\hash.CA1.S0.X[16] ),
    .Q(\hash.CA2.a_dash[16] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[17]$_DFF_P_  (.D(\hash.CA1.S0.X[17] ),
    .Q(\hash.CA2.a_dash[17] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[18]$_DFF_P_  (.D(\hash.CA1.S0.X[18] ),
    .Q(\hash.CA2.a_dash[18] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[19]$_DFF_P_  (.D(\hash.CA1.S0.X[19] ),
    .Q(\hash.CA2.a_dash[19] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[1]$_DFF_P_  (.D(\hash.CA1.S0.X[1] ),
    .Q(\hash.CA2.a_dash[1] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[20]$_DFF_P_  (.D(_06148_),
    .Q(\hash.CA2.a_dash[20] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[21]$_DFF_P_  (.D(_06156_),
    .Q(\hash.CA2.a_dash[21] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[22]$_DFF_P_  (.D(\hash.CA1.S0.X[22] ),
    .Q(\hash.CA2.a_dash[22] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[23]$_DFF_P_  (.D(\hash.CA1.S0.X[23] ),
    .Q(\hash.CA2.a_dash[23] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[24]$_DFF_P_  (.D(_06179_),
    .Q(\hash.CA2.a_dash[24] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[25]$_DFF_P_  (.D(\hash.CA1.S0.X[25] ),
    .Q(\hash.CA2.a_dash[25] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[26]$_DFF_P_  (.D(_06201_),
    .Q(\hash.CA2.a_dash[26] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[27]$_DFF_P_  (.D(_06211_),
    .Q(\hash.CA2.a_dash[27] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[28]$_DFF_P_  (.D(\hash.CA1.S0.X[28] ),
    .Q(\hash.CA2.a_dash[28] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[29]$_DFF_P_  (.D(\hash.CA1.S0.X[29] ),
    .Q(\hash.CA2.a_dash[29] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[2]$_DFF_P_  (.D(\hash.CA1.S0.X[2] ),
    .Q(\hash.CA2.a_dash[2] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[30]$_DFF_P_  (.D(_06234_),
    .Q(\hash.CA2.a_dash[30] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[31]$_DFF_P_  (.D(\hash.CA1.S0.X[31] ),
    .Q(\hash.CA2.a_dash[31] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[3]$_DFF_P_  (.D(\hash.CA1.S0.X[3] ),
    .Q(\hash.CA2.a_dash[3] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[4]$_DFF_P_  (.D(_06010_),
    .Q(\hash.CA2.a_dash[4] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[5]$_DFF_P_  (.D(\hash.CA1.S0.X[5] ),
    .Q(\hash.CA2.a_dash[5] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[6]$_DFF_P_  (.D(\hash.CA1.S0.X[6] ),
    .Q(\hash.CA2.a_dash[6] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[7]$_DFF_P_  (.D(\hash.CA1.S0.X[7] ),
    .Q(\hash.CA2.a_dash[7] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[8]$_DFF_P_  (.D(_06043_),
    .Q(\hash.CA2.a_dash[8] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.a_cap[9]$_DFF_P_  (.D(\hash.CA1.S0.X[9] ),
    .Q(\hash.CA2.a_dash[9] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[0]$_DFF_P_  (.D(\hash.CA1.b[0] ),
    .Q(\hash.CA2.b_dash[0] ),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[10]$_DFF_P_  (.D(\hash.CA1.b[10] ),
    .Q(\hash.CA2.b_dash[10] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[11]$_DFF_P_  (.D(\hash.CA1.b[11] ),
    .Q(\hash.CA2.b_dash[11] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[12]$_DFF_P_  (.D(_06283_),
    .Q(\hash.CA2.b_dash[12] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[13]$_DFF_P_  (.D(\hash.CA1.b[13] ),
    .Q(\hash.CA2.b_dash[13] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[14]$_DFF_P_  (.D(\hash.CA1.b[14] ),
    .Q(\hash.CA2.b_dash[14] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[15]$_DFF_P_  (.D(\hash.CA1.b[15] ),
    .Q(\hash.CA2.b_dash[15] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[16]$_DFF_P_  (.D(\hash.CA1.b[16] ),
    .Q(\hash.CA2.b_dash[16] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[17]$_DFF_P_  (.D(\hash.CA1.b[17] ),
    .Q(\hash.CA2.b_dash[17] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[18]$_DFF_P_  (.D(\hash.CA1.b[18] ),
    .Q(\hash.CA2.b_dash[18] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[19]$_DFF_P_  (.D(_06284_),
    .Q(\hash.CA2.b_dash[19] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[1]$_DFF_P_  (.D(\hash.CA1.b[1] ),
    .Q(\hash.CA2.b_dash[1] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[20]$_DFF_P_  (.D(\hash.CA1.b[20] ),
    .Q(\hash.CA2.b_dash[20] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[21]$_DFF_P_  (.D(\hash.CA1.b[21] ),
    .Q(\hash.CA2.b_dash[21] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[22]$_DFF_P_  (.D(\hash.CA1.b[22] ),
    .Q(\hash.CA2.b_dash[22] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[23]$_DFF_P_  (.D(_06285_),
    .Q(\hash.CA2.b_dash[23] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[24]$_DFF_P_  (.D(\hash.CA1.b[24] ),
    .Q(\hash.CA2.b_dash[24] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[25]$_DFF_P_  (.D(\hash.CA1.b[25] ),
    .Q(\hash.CA2.b_dash[25] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[26]$_DFF_P_  (.D(\hash.CA1.b[26] ),
    .Q(\hash.CA2.b_dash[26] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[27]$_DFF_P_  (.D(\hash.CA1.b[27] ),
    .Q(\hash.CA2.b_dash[27] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[28]$_DFF_P_  (.D(\hash.CA1.b[28] ),
    .Q(\hash.CA2.b_dash[28] ),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[29]$_DFF_P_  (.D(\hash.CA1.b[29] ),
    .Q(\hash.CA2.b_dash[29] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[2]$_DFF_P_  (.D(\hash.CA1.b[2] ),
    .Q(\hash.CA2.b_dash[2] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[30]$_DFF_P_  (.D(\hash.CA1.b[30] ),
    .Q(\hash.CA2.b_dash[30] ),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[31]$_DFF_P_  (.D(\hash.CA1.b[31] ),
    .Q(\hash.CA2.b_dash[31] ),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[3]$_DFF_P_  (.D(\hash.CA1.b[3] ),
    .Q(\hash.CA2.b_dash[3] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[4]$_DFF_P_  (.D(\hash.CA1.b[4] ),
    .Q(\hash.CA2.b_dash[4] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[5]$_DFF_P_  (.D(\hash.CA1.b[5] ),
    .Q(\hash.CA2.b_dash[5] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[6]$_DFF_P_  (.D(\hash.CA1.b[6] ),
    .Q(\hash.CA2.b_dash[6] ),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[7]$_DFF_P_  (.D(\hash.CA1.b[7] ),
    .Q(\hash.CA2.b_dash[7] ),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[8]$_DFF_P_  (.D(_06279_),
    .Q(\hash.CA2.b_dash[8] ),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.b_cap[9]$_DFF_P_  (.D(_06280_),
    .Q(\hash.CA2.b_dash[9] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[0]$_DFF_P_  (.D(\hash.CA1.S1.X[0] ),
    .Q(\hash.CA2.e_dash[0] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[10]$_DFF_P_  (.D(\hash.CA1.S1.X[10] ),
    .Q(\hash.CA2.e_dash[10] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[11]$_DFF_P_  (.D(_06575_),
    .Q(\hash.CA2.e_dash[11] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[12]$_DFF_P_  (.D(\hash.CA1.S1.X[12] ),
    .Q(\hash.CA2.e_dash[12] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[13]$_DFF_P_  (.D(\hash.CA1.S1.X[13] ),
    .Q(\hash.CA2.e_dash[13] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[14]$_DFF_P_  (.D(\hash.CA1.S1.X[14] ),
    .Q(\hash.CA2.e_dash[14] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[15]$_DFF_P_  (.D(_06610_),
    .Q(\hash.CA2.e_dash[15] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[16]$_DFF_P_  (.D(\hash.CA1.S1.X[16] ),
    .Q(\hash.CA2.e_dash[16] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[17]$_DFF_P_  (.D(\hash.CA1.S1.X[17] ),
    .Q(\hash.CA2.e_dash[17] ),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[18]$_DFF_P_  (.D(\hash.CA1.S1.X[18] ),
    .Q(\hash.CA2.e_dash[18] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[19]$_DFF_P_  (.D(\hash.CA1.S1.X[19] ),
    .Q(\hash.CA2.e_dash[19] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.e_cap[1]$_DFF_P_  (.D(\hash.CA1.S1.X[1] ),
    .Q(\hash.CA2.e_dash[1] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[20]$_DFF_P_  (.D(\hash.CA1.S1.X[20] ),
    .Q(\hash.CA2.e_dash[20] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[21]$_DFF_P_  (.D(\hash.CA1.S1.X[21] ),
    .Q(\hash.CA2.e_dash[21] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[22]$_DFF_P_  (.D(\hash.CA1.S1.X[22] ),
    .Q(\hash.CA2.e_dash[22] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[23]$_DFF_P_  (.D(\hash.CA1.S1.X[23] ),
    .Q(\hash.CA2.e_dash[23] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[24]$_DFF_P_  (.D(\hash.CA1.S1.X[24] ),
    .Q(\hash.CA2.e_dash[24] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[25]$_DFF_P_  (.D(net1054),
    .Q(\hash.CA2.e_dash[25] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[26]$_DFF_P_  (.D(_06689_),
    .Q(\hash.CA2.e_dash[26] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[27]$_DFF_P_  (.D(net1124),
    .Q(\hash.CA2.e_dash[27] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[28]$_DFF_P_  (.D(net1097),
    .Q(\hash.CA2.e_dash[28] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[29]$_DFF_P_  (.D(\hash.CA1.S1.X[29] ),
    .Q(\hash.CA2.e_dash[29] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[2]$_DFF_P_  (.D(\hash.CA1.S1.X[2] ),
    .Q(\hash.CA2.e_dash[2] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[30]$_DFF_P_  (.D(net1040),
    .Q(\hash.CA2.e_dash[30] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[31]$_DFF_P_  (.D(\hash.CA1.S1.X[31] ),
    .Q(\hash.CA2.e_dash[31] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.e_cap[3]$_DFF_P_  (.D(\hash.CA1.S1.X[3] ),
    .Q(\hash.CA2.e_dash[3] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[4]$_DFF_P_  (.D(\hash.CA1.S1.X[4] ),
    .Q(\hash.CA2.e_dash[4] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[5]$_DFF_P_  (.D(\hash.CA1.S1.X[5] ),
    .Q(\hash.CA2.e_dash[5] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[6]$_DFF_P_  (.D(\hash.CA1.S1.X[6] ),
    .Q(\hash.CA2.e_dash[6] ),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[7]$_DFF_P_  (.D(\hash.CA1.S1.X[7] ),
    .Q(\hash.CA2.e_dash[7] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[8]$_DFF_P_  (.D(_06552_),
    .Q(\hash.CA2.e_dash[8] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.e_cap[9]$_DFF_P_  (.D(\hash.CA1.S1.X[9] ),
    .Q(\hash.CA2.e_dash[9] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[0]$_DFF_P_  (.D(\hash.CA1.f[0] ),
    .Q(\hash.CA2.f_dash[0] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[10]$_DFF_P_  (.D(\hash.CA1.f[10] ),
    .Q(\hash.CA2.f_dash[10] ),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[11]$_DFF_P_  (.D(\hash.CA1.f[11] ),
    .Q(\hash.CA2.f_dash[11] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[12]$_DFF_P_  (.D(\hash.CA1.f[12] ),
    .Q(\hash.CA2.f_dash[12] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[13]$_DFF_P_  (.D(\hash.CA1.f[13] ),
    .Q(\hash.CA2.f_dash[13] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[14]$_DFF_P_  (.D(\hash.CA1.f[14] ),
    .Q(\hash.CA2.f_dash[14] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[15]$_DFF_P_  (.D(\hash.CA1.f[15] ),
    .Q(\hash.CA2.f_dash[15] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[16]$_DFF_P_  (.D(\hash.CA1.f[16] ),
    .Q(\hash.CA2.f_dash[16] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[17]$_DFF_P_  (.D(\hash.CA1.f[17] ),
    .Q(\hash.CA2.f_dash[17] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[18]$_DFF_P_  (.D(_06467_),
    .Q(\hash.CA2.f_dash[18] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[19]$_DFF_P_  (.D(\hash.CA1.f[19] ),
    .Q(\hash.CA2.f_dash[19] ),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[1]$_DFF_P_  (.D(\hash.CA1.f[1] ),
    .Q(\hash.CA2.f_dash[1] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[20]$_DFF_P_  (.D(\hash.CA1.f[20] ),
    .Q(\hash.CA2.f_dash[20] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[21]$_DFF_P_  (.D(\hash.CA1.f[21] ),
    .Q(\hash.CA2.f_dash[21] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[22]$_DFF_P_  (.D(\hash.CA1.f[22] ),
    .Q(\hash.CA2.f_dash[22] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[23]$_DFF_P_  (.D(\hash.CA1.f[23] ),
    .Q(\hash.CA2.f_dash[23] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[24]$_DFF_P_  (.D(_06487_),
    .Q(\hash.CA2.f_dash[24] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[25]$_DFF_P_  (.D(\hash.CA1.f[25] ),
    .Q(\hash.CA2.f_dash[25] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[26]$_DFF_P_  (.D(\hash.CA1.f[26] ),
    .Q(\hash.CA2.f_dash[26] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[27]$_DFF_P_  (.D(\hash.CA1.f[27] ),
    .Q(\hash.CA2.f_dash[27] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[28]$_DFF_P_  (.D(\hash.CA1.f[28] ),
    .Q(\hash.CA2.f_dash[28] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[29]$_DFF_P_  (.D(\hash.CA1.f[29] ),
    .Q(\hash.CA2.f_dash[29] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[2]$_DFF_P_  (.D(\hash.CA1.f[2] ),
    .Q(\hash.CA2.f_dash[2] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[30]$_DFF_P_  (.D(\hash.CA1.f[30] ),
    .Q(\hash.CA2.f_dash[30] ),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[31]$_DFF_P_  (.D(\hash.CA1.f[31] ),
    .Q(\hash.CA2.f_dash[31] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[3]$_DFF_P_  (.D(\hash.CA1.f[3] ),
    .Q(\hash.CA2.f_dash[3] ),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[4]$_DFF_P_  (.D(\hash.CA1.f[4] ),
    .Q(\hash.CA2.f_dash[4] ),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[5]$_DFF_P_  (.D(\hash.CA1.f[5] ),
    .Q(\hash.CA2.f_dash[5] ),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[6]$_DFF_P_  (.D(\hash.CA1.f[6] ),
    .Q(\hash.CA2.f_dash[6] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[7]$_DFF_P_  (.D(\hash.CA1.f[7] ),
    .Q(\hash.CA2.f_dash[7] ),
    .CLK(clknet_leaf_170_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[8]$_DFF_P_  (.D(\hash.CA1.f[8] ),
    .Q(\hash.CA2.f_dash[8] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.f_cap[9]$_DFF_P_  (.D(_06438_),
    .Q(\hash.CA2.f_dash[9] ),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[0]$_DFFE_PN_  (.D(_00658_),
    .DE(_00906_),
    .Q(net919),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[10]$_DFFE_PN_  (.D(_00659_),
    .DE(_00906_),
    .Q(net930),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[11]$_DFFE_PN_  (.D(_00660_),
    .DE(_00906_),
    .Q(net931),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[12]$_DFFE_PN_  (.D(_00661_),
    .DE(_00906_),
    .Q(net932),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[13]$_DFFE_PN_  (.D(_00662_),
    .DE(_00906_),
    .Q(net933),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[14]$_DFFE_PN_  (.D(_00663_),
    .DE(_00906_),
    .Q(net934),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[15]$_DFFE_PN_  (.D(_00664_),
    .DE(_00906_),
    .Q(net935),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[16]$_DFFE_PN_  (.D(_00665_),
    .DE(_00906_),
    .Q(net937),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[17]$_DFFE_PN_  (.D(_00666_),
    .DE(_00906_),
    .Q(net938),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[18]$_DFFE_PN_  (.D(_00667_),
    .DE(_00906_),
    .Q(net939),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[19]$_DFFE_PN_  (.D(_00668_),
    .DE(_00906_),
    .Q(net940),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[1]$_DFFE_PN_  (.D(_00669_),
    .DE(_00906_),
    .Q(net920),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[20]$_DFFE_PN_  (.D(_00670_),
    .DE(_00906_),
    .Q(net941),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[21]$_DFFE_PN_  (.D(_00671_),
    .DE(_00906_),
    .Q(net942),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[22]$_DFFE_PN_  (.D(_00672_),
    .DE(_00906_),
    .Q(net943),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[23]$_DFFE_PN_  (.D(_00673_),
    .DE(_00906_),
    .Q(net944),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[24]$_DFFE_PN_  (.D(_00674_),
    .DE(_00906_),
    .Q(net945),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[25]$_DFFE_PN_  (.D(_00675_),
    .DE(_00906_),
    .Q(net946),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[26]$_DFFE_PN_  (.D(_00676_),
    .DE(_00906_),
    .Q(net948),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[27]$_DFFE_PN_  (.D(_00677_),
    .DE(_00906_),
    .Q(net949),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[28]$_DFFE_PN_  (.D(_00678_),
    .DE(_00906_),
    .Q(net950),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[29]$_DFFE_PN_  (.D(_00679_),
    .DE(_00906_),
    .Q(net951),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[2]$_DFFE_PN_  (.D(_00680_),
    .DE(_00906_),
    .Q(net921),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[30]$_DFFE_PN_  (.D(_00681_),
    .DE(_00906_),
    .Q(net952),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[31]$_DFFE_PN_  (.D(_00682_),
    .DE(_00906_),
    .Q(net953),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[3]$_DFFE_PN_  (.D(_00683_),
    .DE(_00906_),
    .Q(net922),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[4]$_DFFE_PN_  (.D(_00684_),
    .DE(_00906_),
    .Q(net923),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[5]$_DFFE_PN_  (.D(_00685_),
    .DE(_00906_),
    .Q(net924),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[6]$_DFFE_PN_  (.D(_00686_),
    .DE(_00906_),
    .Q(net926),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[7]$_DFFE_PN_  (.D(_00687_),
    .DE(_00906_),
    .Q(net927),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[8]$_DFFE_PN_  (.D(_00688_),
    .DE(_00906_),
    .Q(net928),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h0_out[9]$_DFFE_PN_  (.D(_00689_),
    .DE(_00906_),
    .Q(net929),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[0]$_DFFE_PN_  (.D(_00690_),
    .DE(_00906_),
    .Q(net883),
    .CLK(clknet_leaf_211_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[10]$_DFFE_PN_  (.D(_00691_),
    .DE(_00906_),
    .Q(net895),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[11]$_DFFE_PN_  (.D(_00692_),
    .DE(_00906_),
    .Q(net896),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[12]$_DFFE_PN_  (.D(_00693_),
    .DE(_00906_),
    .Q(net897),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[13]$_DFFE_PN_  (.D(_00694_),
    .DE(_00906_),
    .Q(net898),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[14]$_DFFE_PN_  (.D(_00695_),
    .DE(_00906_),
    .Q(net899),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[15]$_DFFE_PN_  (.D(_00696_),
    .DE(_00906_),
    .Q(net900),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[16]$_DFFE_PN_  (.D(_00697_),
    .DE(_00906_),
    .Q(net901),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[17]$_DFFE_PN_  (.D(_00698_),
    .DE(_00906_),
    .Q(net902),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[18]$_DFFE_PN_  (.D(_00699_),
    .DE(_00906_),
    .Q(net904),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[19]$_DFFE_PN_  (.D(_00700_),
    .DE(_00906_),
    .Q(net905),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[1]$_DFFE_PN_  (.D(_11575_),
    .DE(_00906_),
    .Q(net884),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[20]$_DFFE_PN_  (.D(_00701_),
    .DE(_00906_),
    .Q(net906),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[21]$_DFFE_PN_  (.D(_00702_),
    .DE(_00906_),
    .Q(net907),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[22]$_DFFE_PN_  (.D(_00703_),
    .DE(_00906_),
    .Q(net908),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[23]$_DFFE_PN_  (.D(_00704_),
    .DE(_00906_),
    .Q(net909),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[24]$_DFFE_PN_  (.D(_00705_),
    .DE(_00906_),
    .Q(net910),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[25]$_DFFE_PN_  (.D(_00706_),
    .DE(_00906_),
    .Q(net911),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[26]$_DFFE_PN_  (.D(_00707_),
    .DE(_00906_),
    .Q(net912),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[27]$_DFFE_PN_  (.D(_00708_),
    .DE(_00906_),
    .Q(net913),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[28]$_DFFE_PN_  (.D(_00709_),
    .DE(_00906_),
    .Q(net915),
    .CLK(clknet_leaf_204_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[29]$_DFFE_PN_  (.D(_00710_),
    .DE(_00906_),
    .Q(net916),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[2]$_DFFE_PN_  (.D(_00711_),
    .DE(_00906_),
    .Q(net885),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[30]$_DFFE_PN_  (.D(_00712_),
    .DE(_00906_),
    .Q(net917),
    .CLK(clknet_leaf_198_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[31]$_DFFE_PN_  (.D(_00713_),
    .DE(_00906_),
    .Q(net918),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[3]$_DFFE_PN_  (.D(_00714_),
    .DE(_00906_),
    .Q(net886),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[4]$_DFFE_PN_  (.D(_00715_),
    .DE(_00906_),
    .Q(net887),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[5]$_DFFE_PN_  (.D(_00716_),
    .DE(_00906_),
    .Q(net888),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[6]$_DFFE_PN_  (.D(_00717_),
    .DE(_00906_),
    .Q(net889),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[7]$_DFFE_PN_  (.D(_00718_),
    .DE(_00906_),
    .Q(net890),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[8]$_DFFE_PN_  (.D(_00719_),
    .DE(_00906_),
    .Q(net893),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h1_out[9]$_DFFE_PN_  (.D(_00720_),
    .DE(_00906_),
    .Q(net894),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[0]$_DFFE_PN_  (.D(\hash.CA1.c[0] ),
    .DE(_00906_),
    .Q(net848),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[10]$_DFFE_PN_  (.D(_00750_),
    .DE(_00906_),
    .Q(net859),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[11]$_DFFE_PN_  (.D(_00722_),
    .DE(_00906_),
    .Q(net860),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[12]$_DFFE_PN_  (.D(_00723_),
    .DE(_00906_),
    .Q(net861),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[13]$_DFFE_PN_  (.D(_00724_),
    .DE(_00906_),
    .Q(net862),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[14]$_DFFE_PN_  (.D(_00725_),
    .DE(_00906_),
    .Q(net863),
    .CLK(clknet_leaf_206_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[15]$_DFFE_PN_  (.D(_00726_),
    .DE(_00906_),
    .Q(net864),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[16]$_DFFE_PN_  (.D(_00727_),
    .DE(_00906_),
    .Q(net865),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[17]$_DFFE_PN_  (.D(_00728_),
    .DE(_00906_),
    .Q(net866),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[18]$_DFFE_PN_  (.D(_00729_),
    .DE(_00906_),
    .Q(net867),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[19]$_DFFE_PN_  (.D(_00730_),
    .DE(_00906_),
    .Q(net868),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[1]$_DFFE_PN_  (.D(_00721_),
    .DE(_00906_),
    .Q(net849),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[20]$_DFFE_PN_  (.D(_00731_),
    .DE(_00906_),
    .Q(net870),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[21]$_DFFE_PN_  (.D(_00732_),
    .DE(_00906_),
    .Q(net871),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[22]$_DFFE_PN_  (.D(_00733_),
    .DE(_00906_),
    .Q(net872),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[23]$_DFFE_PN_  (.D(_00734_),
    .DE(_00906_),
    .Q(net873),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[24]$_DFFE_PN_  (.D(_00735_),
    .DE(_00906_),
    .Q(net874),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[25]$_DFFE_PN_  (.D(_00736_),
    .DE(_00906_),
    .Q(net875),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[26]$_DFFE_PN_  (.D(_00737_),
    .DE(_00906_),
    .Q(net876),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[27]$_DFFE_PN_  (.D(_00738_),
    .DE(_00906_),
    .Q(net877),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[28]$_DFFE_PN_  (.D(_00739_),
    .DE(_00906_),
    .Q(net878),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[29]$_DFFE_PN_  (.D(_00740_),
    .DE(_00906_),
    .Q(net879),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[2]$_DFFE_PN_  (.D(_11576_),
    .DE(_00906_),
    .Q(net850),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[30]$_DFFE_PN_  (.D(_00741_),
    .DE(_00906_),
    .Q(net881),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[31]$_DFFE_PN_  (.D(_00743_),
    .DE(_00906_),
    .Q(net882),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[3]$_DFFE_PN_  (.D(_00742_),
    .DE(_00906_),
    .Q(net851),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[4]$_DFFE_PN_  (.D(_00744_),
    .DE(_00906_),
    .Q(net852),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[5]$_DFFE_PN_  (.D(_00745_),
    .DE(_00906_),
    .Q(net853),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[6]$_DFFE_PN_  (.D(_00746_),
    .DE(_00906_),
    .Q(net854),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[7]$_DFFE_PN_  (.D(_00747_),
    .DE(_00906_),
    .Q(net855),
    .CLK(clknet_leaf_209_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[8]$_DFFE_PN_  (.D(_00748_),
    .DE(_00906_),
    .Q(net856),
    .CLK(clknet_leaf_210_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h2_out[9]$_DFFE_PN_  (.D(_00749_),
    .DE(_00906_),
    .Q(net857),
    .CLK(clknet_leaf_208_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[0]$_DFFE_PN_  (.D(\hash.CA1.d[0] ),
    .DE(_00906_),
    .Q(net812),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[10]$_DFFE_PN_  (.D(_00780_),
    .DE(_00906_),
    .Q(net823),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[11]$_DFFE_PN_  (.D(_00752_),
    .DE(_00906_),
    .Q(net824),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[12]$_DFFE_PN_  (.D(_00753_),
    .DE(_00906_),
    .Q(net826),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[13]$_DFFE_PN_  (.D(_00754_),
    .DE(_00906_),
    .Q(net827),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[14]$_DFFE_PN_  (.D(_00755_),
    .DE(_00906_),
    .Q(net828),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[15]$_DFFE_PN_  (.D(_00756_),
    .DE(_00906_),
    .Q(net829),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[16]$_DFFE_PN_  (.D(_00757_),
    .DE(_00906_),
    .Q(net830),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[17]$_DFFE_PN_  (.D(_00758_),
    .DE(_00906_),
    .Q(net831),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[18]$_DFFE_PN_  (.D(_00759_),
    .DE(_00906_),
    .Q(net832),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[19]$_DFFE_PN_  (.D(_00760_),
    .DE(_00906_),
    .Q(net833),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[1]$_DFFE_PN_  (.D(_00751_),
    .DE(_00906_),
    .Q(net813),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[20]$_DFFE_PN_  (.D(_00761_),
    .DE(_00906_),
    .Q(net834),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[21]$_DFFE_PN_  (.D(_00762_),
    .DE(_00906_),
    .Q(net835),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[22]$_DFFE_PN_  (.D(_00763_),
    .DE(_00906_),
    .Q(net837),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[23]$_DFFE_PN_  (.D(_00764_),
    .DE(_00906_),
    .Q(net838),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[24]$_DFFE_PN_  (.D(_00765_),
    .DE(_00906_),
    .Q(net839),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[25]$_DFFE_PN_  (.D(_00766_),
    .DE(_00906_),
    .Q(net840),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[26]$_DFFE_PN_  (.D(_00767_),
    .DE(_00906_),
    .Q(net841),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[27]$_DFFE_PN_  (.D(_00768_),
    .DE(_00906_),
    .Q(net842),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[28]$_DFFE_PN_  (.D(_00769_),
    .DE(_00906_),
    .Q(net843),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[29]$_DFFE_PN_  (.D(_00770_),
    .DE(_00906_),
    .Q(net844),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[2]$_DFFE_PN_  (.D(_11577_),
    .DE(_00906_),
    .Q(net815),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[30]$_DFFE_PN_  (.D(_00771_),
    .DE(_00906_),
    .Q(net845),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[31]$_DFFE_PN_  (.D(_00773_),
    .DE(_00906_),
    .Q(net846),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[3]$_DFFE_PN_  (.D(_00772_),
    .DE(_00906_),
    .Q(net816),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[4]$_DFFE_PN_  (.D(_00774_),
    .DE(_00906_),
    .Q(net817),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[5]$_DFFE_PN_  (.D(_00775_),
    .DE(_00906_),
    .Q(net818),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[6]$_DFFE_PN_  (.D(_00776_),
    .DE(_00906_),
    .Q(net819),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[7]$_DFFE_PN_  (.D(_00777_),
    .DE(_00906_),
    .Q(net820),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[8]$_DFFE_PN_  (.D(_00778_),
    .DE(_00906_),
    .Q(net821),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h3_out[9]$_DFFE_PN_  (.D(_00779_),
    .DE(_00906_),
    .Q(net822),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[0]$_DFFE_PN_  (.D(_00781_),
    .DE(_00906_),
    .Q(net1032),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[10]$_DFFE_PN_  (.D(_00782_),
    .DE(_00906_),
    .Q(net788),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[11]$_DFFE_PN_  (.D(_00783_),
    .DE(_00906_),
    .Q(net789),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[12]$_DFFE_PN_  (.D(_00784_),
    .DE(_00906_),
    .Q(net790),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[13]$_DFFE_PN_  (.D(_00785_),
    .DE(_00906_),
    .Q(net791),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[14]$_DFFE_PN_  (.D(_00786_),
    .DE(_00906_),
    .Q(net793),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[15]$_DFFE_PN_  (.D(_00787_),
    .DE(_00906_),
    .Q(net794),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[16]$_DFFE_PN_  (.D(_00788_),
    .DE(_00906_),
    .Q(net795),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[17]$_DFFE_PN_  (.D(_00789_),
    .DE(_00906_),
    .Q(net796),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[18]$_DFFE_PN_  (.D(_00790_),
    .DE(_00906_),
    .Q(net797),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[19]$_DFFE_PN_  (.D(_00791_),
    .DE(_00906_),
    .Q(net798),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[1]$_DFFE_PN_  (.D(_00792_),
    .DE(_00906_),
    .Q(net1033),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[20]$_DFFE_PN_  (.D(_00793_),
    .DE(_00906_),
    .Q(net799),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[21]$_DFFE_PN_  (.D(_00794_),
    .DE(_00906_),
    .Q(net800),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[22]$_DFFE_PN_  (.D(_00795_),
    .DE(_00906_),
    .Q(net801),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[23]$_DFFE_PN_  (.D(_00796_),
    .DE(_00906_),
    .Q(net802),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[24]$_DFFE_PN_  (.D(_00797_),
    .DE(_00906_),
    .Q(net804),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[25]$_DFFE_PN_  (.D(_00798_),
    .DE(_00906_),
    .Q(net805),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[26]$_DFFE_PN_  (.D(_00799_),
    .DE(_00906_),
    .Q(net806),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[27]$_DFFE_PN_  (.D(_00800_),
    .DE(_00906_),
    .Q(net807),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[28]$_DFFE_PN_  (.D(_00801_),
    .DE(_00906_),
    .Q(net808),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[29]$_DFFE_PN_  (.D(_00802_),
    .DE(_00906_),
    .Q(net809),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[2]$_DFFE_PN_  (.D(_00803_),
    .DE(_00906_),
    .Q(net1034),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[30]$_DFFE_PN_  (.D(_00804_),
    .DE(_00906_),
    .Q(net810),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[31]$_DFFE_PN_  (.D(_00805_),
    .DE(_00906_),
    .Q(net811),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[3]$_DFFE_PN_  (.D(_00806_),
    .DE(_00906_),
    .Q(net1035),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[4]$_DFFE_PN_  (.D(_00807_),
    .DE(_00906_),
    .Q(net782),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[5]$_DFFE_PN_  (.D(_00808_),
    .DE(_00906_),
    .Q(net783),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[6]$_DFFE_PN_  (.D(_00809_),
    .DE(_00906_),
    .Q(net784),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[7]$_DFFE_PN_  (.D(_00810_),
    .DE(_00906_),
    .Q(net785),
    .CLK(clknet_leaf_195_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[8]$_DFFE_PN_  (.D(_00811_),
    .DE(_00906_),
    .Q(net786),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h4_out[9]$_DFFE_PN_  (.D(_00812_),
    .DE(_00906_),
    .Q(net787),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[0]$_DFFE_PN_  (.D(\hash.CA1.f[0] ),
    .DE(_00906_),
    .Q(net997),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[10]$_DFFE_PN_  (.D(_00841_),
    .DE(_00906_),
    .Q(net1008),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[11]$_DFFE_PN_  (.D(_00842_),
    .DE(_00906_),
    .Q(net1009),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[12]$_DFFE_PN_  (.D(_00814_),
    .DE(_00906_),
    .Q(net1010),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[13]$_DFFE_PN_  (.D(_00815_),
    .DE(_00906_),
    .Q(net1011),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[14]$_DFFE_PN_  (.D(_00816_),
    .DE(_00906_),
    .Q(net1012),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[15]$_DFFE_PN_  (.D(_00817_),
    .DE(_00906_),
    .Q(net1013),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[16]$_DFFE_PN_  (.D(_00818_),
    .DE(_00906_),
    .Q(net1015),
    .CLK(clknet_leaf_165_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[17]$_DFFE_PN_  (.D(_00819_),
    .DE(_00906_),
    .Q(net1016),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[18]$_DFFE_PN_  (.D(_00820_),
    .DE(_00906_),
    .Q(net1017),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[19]$_DFFE_PN_  (.D(_00821_),
    .DE(_00906_),
    .Q(net1018),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[1]$_DFFE_PN_  (.D(\hash.CA1.f[1] ),
    .DE(_00906_),
    .Q(net998),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[20]$_DFFE_PN_  (.D(_00822_),
    .DE(_00906_),
    .Q(net1019),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[21]$_DFFE_PN_  (.D(_00823_),
    .DE(_00906_),
    .Q(net1020),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[22]$_DFFE_PN_  (.D(_00825_),
    .DE(_00906_),
    .Q(net1021),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[23]$_DFFE_PN_  (.D(_00826_),
    .DE(_00906_),
    .Q(net1022),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[24]$_DFFE_PN_  (.D(_00827_),
    .DE(_00906_),
    .Q(net1023),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[25]$_DFFE_PN_  (.D(_00828_),
    .DE(_00906_),
    .Q(net1024),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[26]$_DFFE_PN_  (.D(_00829_),
    .DE(_00906_),
    .Q(net1026),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[27]$_DFFE_PN_  (.D(_00830_),
    .DE(_00906_),
    .Q(net1027),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[28]$_DFFE_PN_  (.D(_00831_),
    .DE(_00906_),
    .Q(net1028),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[29]$_DFFE_PN_  (.D(_00832_),
    .DE(_00906_),
    .Q(net1029),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[2]$_DFFE_PN_  (.D(_00813_),
    .DE(_00906_),
    .Q(net999),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[30]$_DFFE_PN_  (.D(_00833_),
    .DE(_00906_),
    .Q(net1030),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[31]$_DFFE_PN_  (.D(_00834_),
    .DE(_00906_),
    .Q(net1031),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[3]$_DFFE_PN_  (.D(_00824_),
    .DE(_00906_),
    .Q(net1000),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[4]$_DFFE_PN_  (.D(_00835_),
    .DE(_00906_),
    .Q(net1001),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[5]$_DFFE_PN_  (.D(_00836_),
    .DE(_00906_),
    .Q(net1002),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[6]$_DFFE_PN_  (.D(_00837_),
    .DE(_00906_),
    .Q(net1004),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[7]$_DFFE_PN_  (.D(_00838_),
    .DE(_00906_),
    .Q(net1005),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[8]$_DFFE_PN_  (.D(_00839_),
    .DE(_00906_),
    .Q(net1006),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h5_out[9]$_DFFE_PN_  (.D(_00840_),
    .DE(_00906_),
    .Q(net1007),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[0]$_DFFE_PN_  (.D(_00843_),
    .DE(_00906_),
    .Q(net962),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[10]$_DFFE_PN_  (.D(_00844_),
    .DE(_00906_),
    .Q(net973),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[11]$_DFFE_PN_  (.D(_00845_),
    .DE(_00906_),
    .Q(net974),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[12]$_DFFE_PN_  (.D(_00846_),
    .DE(_00906_),
    .Q(net975),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[13]$_DFFE_PN_  (.D(_00847_),
    .DE(_00906_),
    .Q(net976),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[14]$_DFFE_PN_  (.D(_00848_),
    .DE(_00906_),
    .Q(net977),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[15]$_DFFE_PN_  (.D(_00849_),
    .DE(_00906_),
    .Q(net978),
    .CLK(clknet_leaf_196_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[16]$_DFFE_PN_  (.D(_00850_),
    .DE(_00906_),
    .Q(net979),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[17]$_DFFE_PN_  (.D(_00851_),
    .DE(_00906_),
    .Q(net980),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[18]$_DFFE_PN_  (.D(_00852_),
    .DE(_00906_),
    .Q(net982),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[19]$_DFFE_PN_  (.D(_00853_),
    .DE(_00906_),
    .Q(net983),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[1]$_DFFE_PN_  (.D(_00854_),
    .DE(_00906_),
    .Q(net963),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[20]$_DFFE_PN_  (.D(_00855_),
    .DE(_00906_),
    .Q(net984),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[21]$_DFFE_PN_  (.D(_00856_),
    .DE(_00906_),
    .Q(net985),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[22]$_DFFE_PN_  (.D(_00857_),
    .DE(_00906_),
    .Q(net986),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[23]$_DFFE_PN_  (.D(_00858_),
    .DE(_00906_),
    .Q(net987),
    .CLK(clknet_leaf_192_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[24]$_DFFE_PN_  (.D(_00859_),
    .DE(_00906_),
    .Q(net988),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[25]$_DFFE_PN_  (.D(_00860_),
    .DE(_00906_),
    .Q(net989),
    .CLK(clknet_leaf_197_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[26]$_DFFE_PN_  (.D(_00861_),
    .DE(_00906_),
    .Q(net990),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[27]$_DFFE_PN_  (.D(_00862_),
    .DE(_00906_),
    .Q(net991),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[28]$_DFFE_PN_  (.D(_00863_),
    .DE(_00906_),
    .Q(net993),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[29]$_DFFE_PN_  (.D(_00864_),
    .DE(_00906_),
    .Q(net994),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[2]$_DFFE_PN_  (.D(_00865_),
    .DE(_00906_),
    .Q(net964),
    .CLK(clknet_leaf_212_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[30]$_DFFE_PN_  (.D(_00866_),
    .DE(_00906_),
    .Q(net995),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[31]$_DFFE_PN_  (.D(_00867_),
    .DE(_00906_),
    .Q(net996),
    .CLK(clknet_leaf_191_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[3]$_DFFE_PN_  (.D(_00868_),
    .DE(_00906_),
    .Q(net965),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[4]$_DFFE_PN_  (.D(_00869_),
    .DE(_00906_),
    .Q(net966),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[5]$_DFFE_PN_  (.D(_00870_),
    .DE(_00906_),
    .Q(net967),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[6]$_DFFE_PN_  (.D(_00871_),
    .DE(_00906_),
    .Q(net968),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[7]$_DFFE_PN_  (.D(_00872_),
    .DE(_00906_),
    .Q(net969),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[8]$_DFFE_PN_  (.D(_00873_),
    .DE(_00906_),
    .Q(net971),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h6_out[9]$_DFFE_PN_  (.D(_00874_),
    .DE(_00906_),
    .Q(net972),
    .CLK(clknet_leaf_194_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[0]$_DFFE_PN_  (.D(_00875_),
    .DE(_00906_),
    .Q(net781),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[10]$_DFFE_PN_  (.D(_00876_),
    .DE(_00906_),
    .Q(net792),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[11]$_DFFE_PN_  (.D(_00877_),
    .DE(_00906_),
    .Q(net803),
    .CLK(clknet_leaf_163_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[12]$_DFFE_PN_  (.D(_00878_),
    .DE(_00906_),
    .Q(net814),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[13]$_DFFE_PN_  (.D(_00879_),
    .DE(_00906_),
    .Q(net825),
    .CLK(clknet_leaf_164_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[14]$_DFFE_PN_  (.D(_00880_),
    .DE(_00906_),
    .Q(net836),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[15]$_DFFE_PN_  (.D(_00881_),
    .DE(_00906_),
    .Q(net847),
    .CLK(clknet_leaf_162_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[16]$_DFFE_PN_  (.D(_00882_),
    .DE(_00906_),
    .Q(net858),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[17]$_DFFE_PN_  (.D(_00883_),
    .DE(_00906_),
    .Q(net869),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[18]$_DFFE_PN_  (.D(_00884_),
    .DE(_00906_),
    .Q(net880),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[19]$_DFFE_PN_  (.D(_00885_),
    .DE(_00906_),
    .Q(net891),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[1]$_DFFE_PN_  (.D(_11578_),
    .DE(_00906_),
    .Q(net892),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[20]$_DFFE_PN_  (.D(_00886_),
    .DE(_00906_),
    .Q(net903),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[21]$_DFFE_PN_  (.D(_00887_),
    .DE(_00906_),
    .Q(net914),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[22]$_DFFE_PN_  (.D(_00888_),
    .DE(_00906_),
    .Q(net925),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[23]$_DFFE_PN_  (.D(_00889_),
    .DE(_00906_),
    .Q(net936),
    .CLK(clknet_leaf_160_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[24]$_DFFE_PN_  (.D(_00890_),
    .DE(_00906_),
    .Q(net947),
    .CLK(clknet_leaf_161_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[25]$_DFFE_PN_  (.D(_00891_),
    .DE(_00906_),
    .Q(net954),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[26]$_DFFE_PN_  (.D(_00892_),
    .DE(_00906_),
    .Q(net955),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[27]$_DFFE_PN_  (.D(_00893_),
    .DE(_00906_),
    .Q(net956),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[28]$_DFFE_PN_  (.D(_00894_),
    .DE(_00906_),
    .Q(net957),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[29]$_DFFE_PN_  (.D(_00895_),
    .DE(_00906_),
    .Q(net958),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[2]$_DFFE_PN_  (.D(_00896_),
    .DE(_00906_),
    .Q(net959),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[30]$_DFFE_PN_  (.D(_00897_),
    .DE(_00906_),
    .Q(net960),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[31]$_DFFE_PN_  (.D(_00898_),
    .DE(_00906_),
    .Q(net961),
    .CLK(clknet_leaf_154_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[3]$_DFFE_PN_  (.D(_00899_),
    .DE(_00906_),
    .Q(net970),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[4]$_DFFE_PN_  (.D(_00900_),
    .DE(_00906_),
    .Q(net981),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[5]$_DFFE_PN_  (.D(_00901_),
    .DE(_00906_),
    .Q(net992),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[6]$_DFFE_PN_  (.D(_00902_),
    .DE(_00906_),
    .Q(net1003),
    .CLK(clknet_leaf_169_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[7]$_DFFE_PN_  (.D(_00903_),
    .DE(_00906_),
    .Q(net1014),
    .CLK(clknet_leaf_168_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[8]$_DFFE_PN_  (.D(_00904_),
    .DE(_00906_),
    .Q(net1025),
    .CLK(clknet_leaf_167_clk));
 sky130_fd_sc_hd__edfxtp_1 \hash.h7_out[9]$_DFFE_PN_  (.D(_00905_),
    .DE(_00906_),
    .Q(net1036),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p1_cap[0]$_DFF_P_  (.D(\hash.CA1.p1[0] ),
    .Q(\hash.CA2.p1[0] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[10]$_DFF_P_  (.D(\hash.CA1.p1[10] ),
    .Q(\hash.CA2.p1[10] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[11]$_DFF_P_  (.D(\hash.CA1.p1[11] ),
    .Q(\hash.CA2.p1[11] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[12]$_DFF_P_  (.D(\hash.CA1.p1[12] ),
    .Q(\hash.CA2.p1[12] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[13]$_DFF_P_  (.D(\hash.CA1.p1[13] ),
    .Q(\hash.CA2.p1[13] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[14]$_DFF_P_  (.D(\hash.CA1.p1[14] ),
    .Q(\hash.CA2.p1[14] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[15]$_DFF_P_  (.D(\hash.CA1.p1[15] ),
    .Q(\hash.CA2.p1[15] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[16]$_DFF_P_  (.D(\hash.CA1.p1[16] ),
    .Q(\hash.CA2.p1[16] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[17]$_DFF_P_  (.D(\hash.CA1.p1[17] ),
    .Q(\hash.CA2.p1[17] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[18]$_DFF_P_  (.D(\hash.CA1.p1[18] ),
    .Q(\hash.CA2.p1[18] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[19]$_DFF_P_  (.D(\hash.CA1.p1[19] ),
    .Q(\hash.CA2.p1[19] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[1]$_DFF_P_  (.D(\hash.CA1.p1[1] ),
    .Q(\hash.CA2.p1[1] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[20]$_DFF_P_  (.D(\hash.CA1.p1[20] ),
    .Q(\hash.CA2.p1[20] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[21]$_DFF_P_  (.D(\hash.CA1.p1[21] ),
    .Q(\hash.CA2.p1[21] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[22]$_DFF_P_  (.D(\hash.CA1.p1[22] ),
    .Q(\hash.CA2.p1[22] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[23]$_DFF_P_  (.D(\hash.CA1.p1[23] ),
    .Q(\hash.CA2.p1[23] ),
    .CLK(clknet_leaf_200_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[24]$_DFF_P_  (.D(\hash.CA1.p1[24] ),
    .Q(\hash.CA2.p1[24] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[25]$_DFF_P_  (.D(\hash.CA1.p1[25] ),
    .Q(\hash.CA2.p1[25] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[26]$_DFF_P_  (.D(\hash.CA1.p1[26] ),
    .Q(\hash.CA2.p1[26] ),
    .CLK(clknet_leaf_207_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[27]$_DFF_P_  (.D(\hash.CA1.p1[27] ),
    .Q(\hash.CA2.p1[27] ),
    .CLK(clknet_leaf_201_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[28]$_DFF_P_  (.D(\hash.CA1.p1[28] ),
    .Q(\hash.CA2.p1[28] ),
    .CLK(clknet_leaf_199_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[29]$_DFF_P_  (.D(\hash.CA1.p1[29] ),
    .Q(\hash.CA2.p1[29] ),
    .CLK(clknet_leaf_202_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[2]$_DFF_P_  (.D(\hash.CA1.p1[2] ),
    .Q(\hash.CA2.p1[2] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[30]$_DFF_P_  (.D(\hash.CA1.p1[30] ),
    .Q(\hash.CA2.p1[30] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[31]$_DFF_P_  (.D(\hash.CA1.p1[31] ),
    .Q(\hash.CA2.p1[31] ),
    .CLK(clknet_leaf_203_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[3]$_DFF_P_  (.D(\hash.CA1.p1[3] ),
    .Q(\hash.CA2.p1[3] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[4]$_DFF_P_  (.D(\hash.CA1.p1[4] ),
    .Q(\hash.CA2.p1[4] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[5]$_DFF_P_  (.D(\hash.CA1.p1[5] ),
    .Q(\hash.CA2.p1[5] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[6]$_DFF_P_  (.D(\hash.CA1.p1[6] ),
    .Q(\hash.CA2.p1[6] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[7]$_DFF_P_  (.D(\hash.CA1.p1[7] ),
    .Q(\hash.CA2.p1[7] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[8]$_DFF_P_  (.D(\hash.CA1.p1[8] ),
    .Q(\hash.CA2.p1[8] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p1_cap[9]$_DFF_P_  (.D(\hash.CA1.p1[9] ),
    .Q(\hash.CA2.p1[9] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[0]$_DFF_P_  (.D(\hash.CA1.p2[0] ),
    .Q(\hash.CA2.S1.X[0] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[10]$_DFF_P_  (.D(\hash.CA1.p2[10] ),
    .Q(\hash.CA2.S1.X[10] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[11]$_DFF_P_  (.D(\hash.CA1.p2[11] ),
    .Q(\hash.CA2.S1.X[11] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[12]$_DFF_P_  (.D(\hash.CA1.p2[12] ),
    .Q(\hash.CA2.S1.X[12] ),
    .CLK(clknet_leaf_173_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[13]$_DFF_P_  (.D(\hash.CA1.p2[13] ),
    .Q(\hash.CA2.S1.X[13] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[14]$_DFF_P_  (.D(\hash.CA1.p2[14] ),
    .Q(\hash.CA2.S1.X[14] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[15]$_DFF_P_  (.D(\hash.CA1.p2[15] ),
    .Q(\hash.CA2.S1.X[15] ),
    .CLK(clknet_leaf_158_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[16]$_DFF_P_  (.D(\hash.CA1.p2[16] ),
    .Q(\hash.CA2.S1.X[16] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[17]$_DFF_P_  (.D(\hash.CA1.p2[17] ),
    .Q(\hash.CA2.S1.X[17] ),
    .CLK(clknet_leaf_174_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p2_cap[18]$_DFF_P_  (.D(\hash.CA1.p2[18] ),
    .Q(\hash.CA2.S1.X[18] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[19]$_DFF_P_  (.D(\hash.CA1.p2[19] ),
    .Q(\hash.CA2.S1.X[19] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[1]$_DFF_P_  (.D(\hash.CA1.p2[1] ),
    .Q(\hash.CA2.S1.X[1] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[20]$_DFF_P_  (.D(\hash.CA1.p2[20] ),
    .Q(\hash.CA2.S1.X[20] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p2_cap[21]$_DFF_P_  (.D(\hash.CA1.p2[21] ),
    .Q(\hash.CA2.S1.X[21] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p2_cap[22]$_DFF_P_  (.D(\hash.CA1.p2[22] ),
    .Q(\hash.CA2.S1.X[22] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p2_cap[23]$_DFF_P_  (.D(\hash.CA1.p2[23] ),
    .Q(\hash.CA2.S1.X[23] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p2_cap[24]$_DFF_P_  (.D(\hash.CA1.p2[24] ),
    .Q(\hash.CA2.S1.X[24] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[25]$_DFF_P_  (.D(\hash.CA1.p2[25] ),
    .Q(\hash.CA2.S1.X[25] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[26]$_DFF_P_  (.D(\hash.CA1.p2[26] ),
    .Q(\hash.CA2.S1.X[26] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[27]$_DFF_P_  (.D(\hash.CA1.p2[27] ),
    .Q(\hash.CA2.S1.X[27] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[28]$_DFF_P_  (.D(\hash.CA1.p2[28] ),
    .Q(\hash.CA2.S1.X[28] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[29]$_DFF_P_  (.D(\hash.CA1.p2[29] ),
    .Q(\hash.CA2.S1.X[29] ),
    .CLK(clknet_leaf_159_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[2]$_DFF_P_  (.D(\hash.CA1.p2[2] ),
    .Q(\hash.CA2.S1.X[2] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[30]$_DFF_P_  (.D(\hash.CA1.p2[30] ),
    .Q(\hash.CA2.S1.X[30] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p2_cap[31]$_DFF_P_  (.D(\hash.CA1.p2[31] ),
    .Q(\hash.CA2.S1.X[31] ),
    .CLK(clknet_leaf_157_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[3]$_DFF_P_  (.D(\hash.CA1.p2[3] ),
    .Q(\hash.CA2.S1.X[3] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[4]$_DFF_P_  (.D(\hash.CA1.p2[4] ),
    .Q(\hash.CA2.S1.X[4] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p2_cap[5]$_DFF_P_  (.D(\hash.CA1.p2[5] ),
    .Q(\hash.CA2.S1.X[5] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[6]$_DFF_P_  (.D(\hash.CA1.p2[6] ),
    .Q(\hash.CA2.S1.X[6] ),
    .CLK(clknet_leaf_172_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[7]$_DFF_P_  (.D(\hash.CA1.p2[7] ),
    .Q(\hash.CA2.S1.X[7] ),
    .CLK(clknet_leaf_166_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[8]$_DFF_P_  (.D(\hash.CA1.p2[8] ),
    .Q(\hash.CA2.S1.X[8] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_4 \hash.p2_cap[9]$_DFF_P_  (.D(\hash.CA1.p2[9] ),
    .Q(\hash.CA2.S1.X[9] ),
    .CLK(clknet_leaf_171_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p3_cap[0]$_DFF_P_  (.D(\hash.CA1.p3[0] ),
    .Q(\hash.CA2.p3[0] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[10]$_DFF_P_  (.D(\hash.CA1.p3[10] ),
    .Q(\hash.CA2.p3[10] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[11]$_DFF_P_  (.D(\hash.CA1.p3[11] ),
    .Q(\hash.CA2.p3[11] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[12]$_DFF_P_  (.D(\hash.CA1.p3[12] ),
    .Q(\hash.CA2.p3[12] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[13]$_DFF_P_  (.D(\hash.CA1.p3[13] ),
    .Q(\hash.CA2.p3[13] ),
    .CLK(clknet_leaf_205_clk));
 sky130_fd_sc_hd__dfxtp_2 \hash.p3_cap[14]$_DFF_P_  (.D(\hash.CA1.p3[14] ),
    .Q(\hash.CA2.p3[14] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[15]$_DFF_P_  (.D(\hash.CA1.p3[15] ),
    .Q(\hash.CA2.p3[15] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[16]$_DFF_P_  (.D(\hash.CA1.p3[16] ),
    .Q(\hash.CA2.p3[16] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[17]$_DFF_P_  (.D(\hash.CA1.p3[17] ),
    .Q(\hash.CA2.p3[17] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[18]$_DFF_P_  (.D(\hash.CA1.p3[18] ),
    .Q(\hash.CA2.p3[18] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[19]$_DFF_P_  (.D(\hash.CA1.p3[19] ),
    .Q(\hash.CA2.p3[19] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[1]$_DFF_P_  (.D(\hash.CA1.p3[1] ),
    .Q(\hash.CA2.p3[1] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[20]$_DFF_P_  (.D(\hash.CA1.p3[20] ),
    .Q(\hash.CA2.p3[20] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[21]$_DFF_P_  (.D(\hash.CA1.p3[21] ),
    .Q(\hash.CA2.p3[21] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[22]$_DFF_P_  (.D(\hash.CA1.p3[22] ),
    .Q(\hash.CA2.p3[22] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[23]$_DFF_P_  (.D(\hash.CA1.p3[23] ),
    .Q(\hash.CA2.p3[23] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[24]$_DFF_P_  (.D(\hash.CA1.p3[24] ),
    .Q(\hash.CA2.p3[24] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[25]$_DFF_P_  (.D(\hash.CA1.p3[25] ),
    .Q(\hash.CA2.p3[25] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[26]$_DFF_P_  (.D(\hash.CA1.p3[26] ),
    .Q(\hash.CA2.p3[26] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[27]$_DFF_P_  (.D(\hash.CA1.p3[27] ),
    .Q(\hash.CA2.p3[27] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[28]$_DFF_P_  (.D(\hash.CA1.p3[28] ),
    .Q(\hash.CA2.p3[28] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[29]$_DFF_P_  (.D(\hash.CA1.p3[29] ),
    .Q(\hash.CA2.p3[29] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[2]$_DFF_P_  (.D(\hash.CA1.p3[2] ),
    .Q(\hash.CA2.p3[2] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[30]$_DFF_P_  (.D(\hash.CA1.p3[30] ),
    .Q(\hash.CA2.p3[30] ),
    .CLK(clknet_leaf_155_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[31]$_DFF_P_  (.D(\hash.CA1.p3[31] ),
    .Q(\hash.CA2.p3[31] ),
    .CLK(clknet_leaf_156_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[3]$_DFF_P_  (.D(\hash.CA1.p3[3] ),
    .Q(\hash.CA2.p3[3] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[4]$_DFF_P_  (.D(\hash.CA1.p3[4] ),
    .Q(\hash.CA2.p3[4] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[5]$_DFF_P_  (.D(\hash.CA1.p3[5] ),
    .Q(\hash.CA2.p3[5] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[6]$_DFF_P_  (.D(\hash.CA1.p3[6] ),
    .Q(\hash.CA2.p3[6] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[7]$_DFF_P_  (.D(\hash.CA1.p3[7] ),
    .Q(\hash.CA2.p3[7] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[8]$_DFF_P_  (.D(\hash.CA1.p3[8] ),
    .Q(\hash.CA2.p3[8] ),
    .CLK(clknet_leaf_219_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p3_cap[9]$_DFF_P_  (.D(\hash.CA1.p3[9] ),
    .Q(\hash.CA2.p3[9] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[0]$_DFF_P_  (.D(\hash.CA1.p4[0] ),
    .Q(\hash.CA2.p4[0] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[10]$_DFF_P_  (.D(\hash.CA1.p4[10] ),
    .Q(\hash.CA2.p4[10] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[11]$_DFF_P_  (.D(\hash.CA1.p4[11] ),
    .Q(\hash.CA2.p4[11] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[12]$_DFF_P_  (.D(\hash.CA1.p4[12] ),
    .Q(\hash.CA2.p4[12] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[13]$_DFF_P_  (.D(\hash.CA1.p4[13] ),
    .Q(\hash.CA2.p4[13] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[14]$_DFF_P_  (.D(\hash.CA1.p4[14] ),
    .Q(\hash.CA2.p4[14] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[15]$_DFF_P_  (.D(\hash.CA1.p4[15] ),
    .Q(\hash.CA2.p4[15] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[16]$_DFF_P_  (.D(\hash.CA1.p4[16] ),
    .Q(\hash.CA2.p4[16] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[17]$_DFF_P_  (.D(\hash.CA1.p4[17] ),
    .Q(\hash.CA2.p4[17] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[18]$_DFF_P_  (.D(\hash.CA1.p4[18] ),
    .Q(\hash.CA2.p4[18] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[19]$_DFF_P_  (.D(\hash.CA1.p4[19] ),
    .Q(\hash.CA2.p4[19] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[1]$_DFF_P_  (.D(\hash.CA1.p4[1] ),
    .Q(\hash.CA2.p4[1] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[20]$_DFF_P_  (.D(\hash.CA1.p4[20] ),
    .Q(\hash.CA2.p4[20] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[21]$_DFF_P_  (.D(\hash.CA1.p4[21] ),
    .Q(\hash.CA2.p4[21] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[22]$_DFF_P_  (.D(\hash.CA1.p4[22] ),
    .Q(\hash.CA2.p4[22] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[23]$_DFF_P_  (.D(\hash.CA1.p4[23] ),
    .Q(\hash.CA2.p4[23] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[24]$_DFF_P_  (.D(\hash.CA1.p4[24] ),
    .Q(\hash.CA2.p4[24] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[25]$_DFF_P_  (.D(\hash.CA1.p4[25] ),
    .Q(\hash.CA2.p4[25] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[26]$_DFF_P_  (.D(\hash.CA1.p4[26] ),
    .Q(\hash.CA2.p4[26] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[27]$_DFF_P_  (.D(\hash.CA1.p4[27] ),
    .Q(\hash.CA2.p4[27] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[28]$_DFF_P_  (.D(\hash.CA1.p4[28] ),
    .Q(\hash.CA2.p4[28] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[29]$_DFF_P_  (.D(\hash.CA1.p4[29] ),
    .Q(\hash.CA2.p4[29] ),
    .CLK(clknet_leaf_188_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[2]$_DFF_P_  (.D(\hash.CA1.p4[2] ),
    .Q(\hash.CA2.p4[2] ),
    .CLK(clknet_leaf_215_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[30]$_DFF_P_  (.D(\hash.CA1.p4[30] ),
    .Q(\hash.CA2.p4[30] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[31]$_DFF_P_  (.D(\hash.CA1.p4[31] ),
    .Q(\hash.CA2.p4[31] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[3]$_DFF_P_  (.D(\hash.CA1.p4[3] ),
    .Q(\hash.CA2.p4[3] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[4]$_DFF_P_  (.D(\hash.CA1.p4[4] ),
    .Q(\hash.CA2.p4[4] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[5]$_DFF_P_  (.D(\hash.CA1.p4[5] ),
    .Q(\hash.CA2.p4[5] ),
    .CLK(clknet_leaf_216_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[6]$_DFF_P_  (.D(\hash.CA1.p4[6] ),
    .Q(\hash.CA2.p4[6] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[7]$_DFF_P_  (.D(\hash.CA1.p4[7] ),
    .Q(\hash.CA2.p4[7] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[8]$_DFF_P_  (.D(\hash.CA1.p4[8] ),
    .Q(\hash.CA2.p4[8] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p4_cap[9]$_DFF_P_  (.D(\hash.CA1.p4[9] ),
    .Q(\hash.CA2.p4[9] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[0]$_DFF_P_  (.D(\hash.CA1.p5[0] ),
    .Q(\hash.CA2.p5[0] ),
    .CLK(clknet_leaf_213_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[10]$_DFF_P_  (.D(\hash.CA1.p5[10] ),
    .Q(\hash.CA2.p5[10] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[11]$_DFF_P_  (.D(\hash.CA1.p5[11] ),
    .Q(\hash.CA2.p5[11] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[12]$_DFF_P_  (.D(\hash.CA1.p5[12] ),
    .Q(\hash.CA2.p5[12] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[13]$_DFF_P_  (.D(\hash.CA1.p5[13] ),
    .Q(\hash.CA2.p5[13] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[14]$_DFF_P_  (.D(\hash.CA1.p5[14] ),
    .Q(\hash.CA2.p5[14] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[15]$_DFF_P_  (.D(\hash.CA1.p5[15] ),
    .Q(\hash.CA2.p5[15] ),
    .CLK(clknet_leaf_187_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[16]$_DFF_P_  (.D(\hash.CA1.p5[16] ),
    .Q(\hash.CA2.p5[16] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[17]$_DFF_P_  (.D(\hash.CA1.p5[17] ),
    .Q(\hash.CA2.p5[17] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[18]$_DFF_P_  (.D(\hash.CA1.p5[18] ),
    .Q(\hash.CA2.p5[18] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[19]$_DFF_P_  (.D(\hash.CA1.p5[19] ),
    .Q(\hash.CA2.p5[19] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[1]$_DFF_P_  (.D(\hash.CA1.p5[1] ),
    .Q(\hash.CA2.p5[1] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[20]$_DFF_P_  (.D(\hash.CA1.p5[20] ),
    .Q(\hash.CA2.p5[20] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[21]$_DFF_P_  (.D(\hash.CA1.p5[21] ),
    .Q(\hash.CA2.p5[21] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[22]$_DFF_P_  (.D(\hash.CA1.p5[22] ),
    .Q(\hash.CA2.p5[22] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[23]$_DFF_P_  (.D(\hash.CA1.p5[23] ),
    .Q(\hash.CA2.p5[23] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[24]$_DFF_P_  (.D(\hash.CA1.p5[24] ),
    .Q(\hash.CA2.p5[24] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[25]$_DFF_P_  (.D(\hash.CA1.p5[25] ),
    .Q(\hash.CA2.p5[25] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[26]$_DFF_P_  (.D(\hash.CA1.p5[26] ),
    .Q(\hash.CA2.p5[26] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[27]$_DFF_P_  (.D(\hash.CA1.p5[27] ),
    .Q(\hash.CA2.p5[27] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[28]$_DFF_P_  (.D(\hash.CA1.p5[28] ),
    .Q(\hash.CA2.p5[28] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[29]$_DFF_P_  (.D(\hash.CA1.p5[29] ),
    .Q(\hash.CA2.p5[29] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[2]$_DFF_P_  (.D(\hash.CA1.p5[2] ),
    .Q(\hash.CA2.p5[2] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[30]$_DFF_P_  (.D(\hash.CA1.p5[30] ),
    .Q(\hash.CA2.p5[30] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[31]$_DFF_P_  (.D(\hash.CA1.p5[31] ),
    .Q(\hash.CA2.p5[31] ),
    .CLK(clknet_leaf_189_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[3]$_DFF_P_  (.D(\hash.CA1.p5[3] ),
    .Q(\hash.CA2.p5[3] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[4]$_DFF_P_  (.D(\hash.CA1.p5[4] ),
    .Q(\hash.CA2.p5[4] ),
    .CLK(clknet_leaf_214_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[5]$_DFF_P_  (.D(\hash.CA1.p5[5] ),
    .Q(\hash.CA2.p5[5] ),
    .CLK(clknet_leaf_190_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[6]$_DFF_P_  (.D(\hash.CA1.p5[6] ),
    .Q(\hash.CA2.p5[6] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[7]$_DFF_P_  (.D(\hash.CA1.p5[7] ),
    .Q(\hash.CA2.p5[7] ),
    .CLK(clknet_leaf_217_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[8]$_DFF_P_  (.D(\hash.CA1.p5[8] ),
    .Q(\hash.CA2.p5[8] ),
    .CLK(clknet_leaf_186_clk));
 sky130_fd_sc_hd__dfxtp_1 \hash.p5_cap[9]$_DFF_P_  (.D(\hash.CA1.p5[9] ),
    .Q(\hash.CA2.p5[9] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[0]$_SDFF_PP0_  (.D(_00969_),
    .Q(\hash.CA1.k_i1[0] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[10]$_SDFF_PP1_  (.D(_00970_),
    .Q(\hash.CA1.k_i1[10] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[11]$_SDFF_PP1_  (.D(_00971_),
    .Q(\hash.CA1.k_i1[11] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[12]$_SDFF_PP0_  (.D(_00972_),
    .Q(\hash.CA1.k_i1[12] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[13]$_SDFF_PP1_  (.D(_00973_),
    .Q(\hash.CA1.k_i1[13] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[14]$_SDFF_PP0_  (.D(_00974_),
    .Q(\hash.CA1.k_i1[14] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[15]$_SDFF_PP0_  (.D(_00975_),
    .Q(\hash.CA1.k_i1[15] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[16]$_SDFF_PP0_  (.D(_00976_),
    .Q(\hash.CA1.k_i1[16] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[17]$_SDFF_PP1_  (.D(_00977_),
    .Q(\hash.CA1.k_i1[17] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[18]$_SDFF_PP0_  (.D(_00978_),
    .Q(\hash.CA1.k_i1[18] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[19]$_SDFF_PP1_  (.D(_00979_),
    .Q(\hash.CA1.k_i1[19] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[1]$_SDFF_PP0_  (.D(_00980_),
    .Q(\hash.CA1.k_i1[1] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[20]$_SDFF_PP0_  (.D(_00981_),
    .Q(\hash.CA1.k_i1[20] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[21]$_SDFF_PP0_  (.D(_00982_),
    .Q(\hash.CA1.k_i1[21] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[22]$_SDFF_PP0_  (.D(_00983_),
    .Q(\hash.CA1.k_i1[22] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[23]$_SDFF_PP1_  (.D(_00984_),
    .Q(\hash.CA1.k_i1[23] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[24]$_SDFF_PP0_  (.D(_00985_),
    .Q(\hash.CA1.k_i1[24] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[25]$_SDFF_PP1_  (.D(_00986_),
    .Q(\hash.CA1.k_i1[25] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[26]$_SDFF_PP0_  (.D(_00987_),
    .Q(\hash.CA1.k_i1[26] ),
    .CLK(clknet_leaf_151_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[27]$_SDFF_PP0_  (.D(_00988_),
    .Q(\hash.CA1.k_i1[27] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[28]$_SDFF_PP0_  (.D(_00989_),
    .Q(\hash.CA1.k_i1[28] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[29]$_SDFF_PP0_  (.D(_00990_),
    .Q(\hash.CA1.k_i1[29] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[2]$_SDFF_PP0_  (.D(_00991_),
    .Q(\hash.CA1.k_i1[2] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[30]$_SDFF_PP1_  (.D(_00992_),
    .Q(\hash.CA1.k_i1[30] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[31]$_SDFF_PP0_  (.D(_00993_),
    .Q(\hash.CA1.k_i1[31] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[3]$_SDFF_PP1_  (.D(_00994_),
    .Q(\hash.CA1.k_i1[3] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[4]$_SDFF_PP1_  (.D(_00995_),
    .Q(\hash.CA1.k_i1[4] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[5]$_SDFF_PP0_  (.D(_00996_),
    .Q(\hash.CA1.k_i1[5] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[6]$_SDFF_PP0_  (.D(_00997_),
    .Q(\hash.CA1.k_i1[6] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[7]$_SDFF_PP1_  (.D(_00998_),
    .Q(\hash.CA1.k_i1[7] ),
    .CLK(clknet_leaf_134_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[8]$_SDFF_PP1_  (.D(_00999_),
    .Q(\hash.CA1.k_i1[8] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value1[9]$_SDFF_PP1_  (.D(_01000_),
    .Q(\hash.CA1.k_i1[9] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[0]$_SDFF_PP1_  (.D(_01001_),
    .Q(\hash.CA1.k_i2[0] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[10]$_SDFF_PP1_  (.D(_01002_),
    .Q(\hash.CA1.k_i2[10] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[11]$_SDFF_PP0_  (.D(_01003_),
    .Q(\hash.CA1.k_i2[11] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[12]$_SDFF_PP0_  (.D(_01004_),
    .Q(\hash.CA1.k_i2[12] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[13]$_SDFF_PP0_  (.D(_01005_),
    .Q(\hash.CA1.k_i2[13] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[14]$_SDFF_PP1_  (.D(_01006_),
    .Q(\hash.CA1.k_i2[14] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[15]$_SDFF_PP0_  (.D(_01007_),
    .Q(\hash.CA1.k_i2[15] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[16]$_SDFF_PP1_  (.D(_01008_),
    .Q(\hash.CA1.k_i2[16] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[17]$_SDFF_PP1_  (.D(_01009_),
    .Q(\hash.CA1.k_i2[17] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[18]$_SDFF_PP1_  (.D(_01010_),
    .Q(\hash.CA1.k_i2[18] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[19]$_SDFF_PP0_  (.D(_01011_),
    .Q(\hash.CA1.k_i2[19] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[1]$_SDFF_PP0_  (.D(_01012_),
    .Q(\hash.CA1.k_i2[1] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[20]$_SDFF_PP1_  (.D(_01013_),
    .Q(\hash.CA1.k_i2[20] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[21]$_SDFF_PP1_  (.D(_01014_),
    .Q(\hash.CA1.k_i2[21] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[22]$_SDFF_PP0_  (.D(_01015_),
    .Q(\hash.CA1.k_i2[22] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[23]$_SDFF_PP0_  (.D(_01016_),
    .Q(\hash.CA1.k_i2[23] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[24]$_SDFF_PP1_  (.D(_01017_),
    .Q(\hash.CA1.k_i2[24] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[25]$_SDFF_PP0_  (.D(_01018_),
    .Q(\hash.CA1.k_i2[25] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[26]$_SDFF_PP0_  (.D(_01019_),
    .Q(\hash.CA1.k_i2[26] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[27]$_SDFF_PP0_  (.D(_01020_),
    .Q(\hash.CA1.k_i2[27] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[28]$_SDFF_PP1_  (.D(_01021_),
    .Q(\hash.CA1.k_i2[28] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[29]$_SDFF_PP1_  (.D(_01022_),
    .Q(\hash.CA1.k_i2[29] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[2]$_SDFF_PP0_  (.D(_01023_),
    .Q(\hash.CA1.k_i2[2] ),
    .CLK(clknet_leaf_218_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[30]$_SDFF_PP1_  (.D(_01024_),
    .Q(\hash.CA1.k_i2[30] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[31]$_SDFF_PP0_  (.D(_01025_),
    .Q(\hash.CA1.k_i2[31] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[3]$_SDFF_PP0_  (.D(_01026_),
    .Q(\hash.CA1.k_i2[3] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[4]$_SDFF_PP1_  (.D(_01027_),
    .Q(\hash.CA1.k_i2[4] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[5]$_SDFF_PP0_  (.D(_01028_),
    .Q(\hash.CA1.k_i2[5] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[6]$_SDFF_PP0_  (.D(_01029_),
    .Q(\hash.CA1.k_i2[6] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[7]$_SDFF_PP1_  (.D(_01030_),
    .Q(\hash.CA1.k_i2[7] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[8]$_SDFF_PP0_  (.D(_01031_),
    .Q(\hash.CA1.k_i2[8] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 \k_value2[9]$_SDFF_PP0_  (.D(_01032_),
    .Q(\hash.CA1.k_i2[9] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \ready$_DFF_P_  (.D(ready_dash),
    .Q(net1037),
    .CLK(clknet_leaf_193_clk));
 sky130_fd_sc_hd__dfxtp_1 \ready_dash$_SDFF_PP0_  (.D(_01033_),
    .Q(ready_dash),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 \reset_hash$_DFF_P_  (.D(net1038),
    .Q(reset_hash),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__dfxtp_1 \reset_hash_dash$_DFF_P_  (.D(net349),
    .Q(\hash.reset ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][0]$_DFFE_PP_  (.D(_00129_),
    .DE(_00127_),
    .Q(\w[0][0] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][10]$_DFFE_PP_  (.D(_00130_),
    .DE(_00127_),
    .Q(\w[0][10] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][11]$_DFFE_PP_  (.D(_00131_),
    .DE(_00127_),
    .Q(\w[0][11] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][12]$_DFFE_PP_  (.D(_00132_),
    .DE(_00127_),
    .Q(\w[0][12] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][13]$_DFFE_PP_  (.D(_00133_),
    .DE(_00127_),
    .Q(\w[0][13] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][14]$_DFFE_PP_  (.D(_00134_),
    .DE(_00127_),
    .Q(\w[0][14] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][15]$_DFFE_PP_  (.D(_00135_),
    .DE(_00127_),
    .Q(\w[0][15] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][16]$_DFFE_PP_  (.D(_00136_),
    .DE(_00127_),
    .Q(\w[0][16] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][17]$_DFFE_PP_  (.D(_00137_),
    .DE(_00127_),
    .Q(\w[0][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][18]$_DFFE_PP_  (.D(_00138_),
    .DE(_00127_),
    .Q(\w[0][18] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][19]$_DFFE_PP_  (.D(_00139_),
    .DE(_00127_),
    .Q(\w[0][19] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][1]$_DFFE_PP_  (.D(_00140_),
    .DE(_00127_),
    .Q(\w[0][1] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][20]$_DFFE_PP_  (.D(_00141_),
    .DE(_00127_),
    .Q(\w[0][20] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][21]$_DFFE_PP_  (.D(_00142_),
    .DE(_00127_),
    .Q(\w[0][21] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][22]$_DFFE_PP_  (.D(_00143_),
    .DE(_00127_),
    .Q(\w[0][22] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][23]$_DFFE_PP_  (.D(_00144_),
    .DE(_00127_),
    .Q(\w[0][23] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][24]$_DFFE_PP_  (.D(_00145_),
    .DE(_00127_),
    .Q(\w[0][24] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][25]$_DFFE_PP_  (.D(_00146_),
    .DE(_00127_),
    .Q(\w[0][25] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][26]$_DFFE_PP_  (.D(_00147_),
    .DE(_00127_),
    .Q(\w[0][26] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][27]$_DFFE_PP_  (.D(_00148_),
    .DE(_00127_),
    .Q(\w[0][27] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][28]$_DFFE_PP_  (.D(_00149_),
    .DE(_00127_),
    .Q(\w[0][28] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][29]$_DFFE_PP_  (.D(_00150_),
    .DE(_00127_),
    .Q(\w[0][29] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][2]$_DFFE_PP_  (.D(_00151_),
    .DE(_00127_),
    .Q(\w[0][2] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][30]$_DFFE_PP_  (.D(_00152_),
    .DE(_00127_),
    .Q(\w[0][30] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][31]$_DFFE_PP_  (.D(_00153_),
    .DE(_00127_),
    .Q(\w[0][31] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][3]$_DFFE_PP_  (.D(_00154_),
    .DE(_00127_),
    .Q(\w[0][3] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][4]$_DFFE_PP_  (.D(_00155_),
    .DE(_00127_),
    .Q(\w[0][4] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][5]$_DFFE_PP_  (.D(_00156_),
    .DE(_00127_),
    .Q(\w[0][5] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][6]$_DFFE_PP_  (.D(_00157_),
    .DE(_00127_),
    .Q(\w[0][6] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][7]$_DFFE_PP_  (.D(_00158_),
    .DE(_00127_),
    .Q(\w[0][7] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][8]$_DFFE_PP_  (.D(_00159_),
    .DE(_00127_),
    .Q(\w[0][8] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[0][9]$_DFFE_PP_  (.D(_00160_),
    .DE(_00127_),
    .Q(\w[0][9] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][0]$_DFFE_PP_  (.D(_00161_),
    .DE(_00126_),
    .Q(\w[10][0] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][10]$_DFFE_PP_  (.D(_00162_),
    .DE(_00126_),
    .Q(\w[10][10] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][11]$_DFFE_PP_  (.D(_00163_),
    .DE(_00126_),
    .Q(\w[10][11] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][12]$_DFFE_PP_  (.D(_00164_),
    .DE(_00126_),
    .Q(\w[10][12] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][13]$_DFFE_PP_  (.D(_00165_),
    .DE(_00126_),
    .Q(\w[10][13] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][14]$_DFFE_PP_  (.D(_00166_),
    .DE(_00126_),
    .Q(\w[10][14] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][15]$_DFFE_PP_  (.D(_00167_),
    .DE(_00126_),
    .Q(\w[10][15] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][16]$_DFFE_PP_  (.D(_00168_),
    .DE(_00126_),
    .Q(\w[10][16] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][17]$_DFFE_PP_  (.D(_00169_),
    .DE(_00126_),
    .Q(\w[10][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][18]$_DFFE_PP_  (.D(_00170_),
    .DE(_00126_),
    .Q(\w[10][18] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][19]$_DFFE_PP_  (.D(_00171_),
    .DE(_00126_),
    .Q(\w[10][19] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][1]$_DFFE_PP_  (.D(_00172_),
    .DE(_00126_),
    .Q(\w[10][1] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][20]$_DFFE_PP_  (.D(_00173_),
    .DE(_00126_),
    .Q(\w[10][20] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][21]$_DFFE_PP_  (.D(_00174_),
    .DE(_00126_),
    .Q(\w[10][21] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][22]$_DFFE_PP_  (.D(_00175_),
    .DE(_00126_),
    .Q(\w[10][22] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][23]$_DFFE_PP_  (.D(_00176_),
    .DE(_00126_),
    .Q(\w[10][23] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][24]$_DFFE_PP_  (.D(_00177_),
    .DE(_00126_),
    .Q(\w[10][24] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][25]$_DFFE_PP_  (.D(_00178_),
    .DE(_00126_),
    .Q(\w[10][25] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][26]$_DFFE_PP_  (.D(_00179_),
    .DE(_00126_),
    .Q(\w[10][26] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][27]$_DFFE_PP_  (.D(_00180_),
    .DE(_00126_),
    .Q(\w[10][27] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][28]$_DFFE_PP_  (.D(_00181_),
    .DE(_00126_),
    .Q(\w[10][28] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][29]$_DFFE_PP_  (.D(_00182_),
    .DE(_00126_),
    .Q(\w[10][29] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][2]$_DFFE_PP_  (.D(_00183_),
    .DE(_00126_),
    .Q(\w[10][2] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][30]$_DFFE_PP_  (.D(_00184_),
    .DE(_00126_),
    .Q(\w[10][30] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][31]$_DFFE_PP_  (.D(_00185_),
    .DE(_00126_),
    .Q(\w[10][31] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][3]$_DFFE_PP_  (.D(_00186_),
    .DE(_00126_),
    .Q(\w[10][3] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][4]$_DFFE_PP_  (.D(_00187_),
    .DE(_00126_),
    .Q(\w[10][4] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][5]$_DFFE_PP_  (.D(_00188_),
    .DE(_00126_),
    .Q(\w[10][5] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][6]$_DFFE_PP_  (.D(_00189_),
    .DE(_00126_),
    .Q(\w[10][6] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][7]$_DFFE_PP_  (.D(_00190_),
    .DE(_00126_),
    .Q(\w[10][7] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][8]$_DFFE_PP_  (.D(_00191_),
    .DE(_00126_),
    .Q(\w[10][8] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[10][9]$_DFFE_PP_  (.D(_00192_),
    .DE(_00126_),
    .Q(\w[10][9] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][0]$_DFFE_PP_  (.D(_00193_),
    .DE(_00095_),
    .Q(\w[11][0] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][10]$_DFFE_PP_  (.D(_00194_),
    .DE(_00095_),
    .Q(\w[11][10] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][11]$_DFFE_PP_  (.D(_00195_),
    .DE(_00095_),
    .Q(\w[11][11] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][12]$_DFFE_PP_  (.D(_00196_),
    .DE(_00095_),
    .Q(\w[11][12] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][13]$_DFFE_PP_  (.D(_00197_),
    .DE(_00095_),
    .Q(\w[11][13] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][14]$_DFFE_PP_  (.D(_00198_),
    .DE(_00095_),
    .Q(\w[11][14] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][15]$_DFFE_PP_  (.D(_00199_),
    .DE(_00095_),
    .Q(\w[11][15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][16]$_DFFE_PP_  (.D(_00200_),
    .DE(_00095_),
    .Q(\w[11][16] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][17]$_DFFE_PP_  (.D(_00201_),
    .DE(_00095_),
    .Q(\w[11][17] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][18]$_DFFE_PP_  (.D(_00202_),
    .DE(_00095_),
    .Q(\w[11][18] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][19]$_DFFE_PP_  (.D(_00203_),
    .DE(_00095_),
    .Q(\w[11][19] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][1]$_DFFE_PP_  (.D(_00204_),
    .DE(_00095_),
    .Q(\w[11][1] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][20]$_DFFE_PP_  (.D(_00205_),
    .DE(_00095_),
    .Q(\w[11][20] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][21]$_DFFE_PP_  (.D(_00206_),
    .DE(_00095_),
    .Q(\w[11][21] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][22]$_DFFE_PP_  (.D(_00207_),
    .DE(_00095_),
    .Q(\w[11][22] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][23]$_DFFE_PP_  (.D(_00208_),
    .DE(_00095_),
    .Q(\w[11][23] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][24]$_DFFE_PP_  (.D(_00209_),
    .DE(_00095_),
    .Q(\w[11][24] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][25]$_DFFE_PP_  (.D(_00210_),
    .DE(_00095_),
    .Q(\w[11][25] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][26]$_DFFE_PP_  (.D(_00211_),
    .DE(_00095_),
    .Q(\w[11][26] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][27]$_DFFE_PP_  (.D(_00212_),
    .DE(_00095_),
    .Q(\w[11][27] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][28]$_DFFE_PP_  (.D(_00213_),
    .DE(_00095_),
    .Q(\w[11][28] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][29]$_DFFE_PP_  (.D(_00214_),
    .DE(_00095_),
    .Q(\w[11][29] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][2]$_DFFE_PP_  (.D(_00215_),
    .DE(_00095_),
    .Q(\w[11][2] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][30]$_DFFE_PP_  (.D(_00216_),
    .DE(_00095_),
    .Q(\w[11][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][31]$_DFFE_PP_  (.D(_00217_),
    .DE(_00095_),
    .Q(\w[11][31] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][3]$_DFFE_PP_  (.D(_00218_),
    .DE(_00095_),
    .Q(\w[11][3] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][4]$_DFFE_PP_  (.D(_00219_),
    .DE(_00095_),
    .Q(\w[11][4] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][5]$_DFFE_PP_  (.D(_00220_),
    .DE(_00095_),
    .Q(\w[11][5] ),
    .CLK(clknet_leaf_290_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][6]$_DFFE_PP_  (.D(_00221_),
    .DE(_00095_),
    .Q(\w[11][6] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][7]$_DFFE_PP_  (.D(_00222_),
    .DE(_00095_),
    .Q(\w[11][7] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][8]$_DFFE_PP_  (.D(_00223_),
    .DE(_00095_),
    .Q(\w[11][8] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[11][9]$_DFFE_PP_  (.D(_00224_),
    .DE(_00095_),
    .Q(\w[11][9] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][0]$_DFFE_PP_  (.D(_00225_),
    .DE(_00125_),
    .Q(\w[12][0] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][10]$_DFFE_PP_  (.D(_00226_),
    .DE(_00125_),
    .Q(\w[12][10] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][11]$_DFFE_PP_  (.D(_00227_),
    .DE(_00125_),
    .Q(\w[12][11] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][12]$_DFFE_PP_  (.D(_00228_),
    .DE(_00125_),
    .Q(\w[12][12] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][13]$_DFFE_PP_  (.D(_00229_),
    .DE(_00125_),
    .Q(\w[12][13] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][14]$_DFFE_PP_  (.D(_00230_),
    .DE(_00125_),
    .Q(\w[12][14] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][15]$_DFFE_PP_  (.D(_00231_),
    .DE(_00125_),
    .Q(\w[12][15] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][16]$_DFFE_PP_  (.D(_00232_),
    .DE(_00125_),
    .Q(\w[12][16] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][17]$_DFFE_PP_  (.D(_00233_),
    .DE(_00125_),
    .Q(\w[12][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][18]$_DFFE_PP_  (.D(_00234_),
    .DE(_00125_),
    .Q(\w[12][18] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][19]$_DFFE_PP_  (.D(_00235_),
    .DE(_00125_),
    .Q(\w[12][19] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][1]$_DFFE_PP_  (.D(_00236_),
    .DE(_00125_),
    .Q(\w[12][1] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][20]$_DFFE_PP_  (.D(_00237_),
    .DE(_00125_),
    .Q(\w[12][20] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][21]$_DFFE_PP_  (.D(_00238_),
    .DE(_00125_),
    .Q(\w[12][21] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][22]$_DFFE_PP_  (.D(_00239_),
    .DE(_00125_),
    .Q(\w[12][22] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][23]$_DFFE_PP_  (.D(_00240_),
    .DE(_00125_),
    .Q(\w[12][23] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][24]$_DFFE_PP_  (.D(_00241_),
    .DE(_00125_),
    .Q(\w[12][24] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][25]$_DFFE_PP_  (.D(_00242_),
    .DE(_00125_),
    .Q(\w[12][25] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][26]$_DFFE_PP_  (.D(_00243_),
    .DE(_00125_),
    .Q(\w[12][26] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][27]$_DFFE_PP_  (.D(_00244_),
    .DE(_00125_),
    .Q(\w[12][27] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][28]$_DFFE_PP_  (.D(_00245_),
    .DE(_00125_),
    .Q(\w[12][28] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][29]$_DFFE_PP_  (.D(_00246_),
    .DE(_00125_),
    .Q(\w[12][29] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][2]$_DFFE_PP_  (.D(_00247_),
    .DE(_00125_),
    .Q(\w[12][2] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][30]$_DFFE_PP_  (.D(_00248_),
    .DE(_00125_),
    .Q(\w[12][30] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][31]$_DFFE_PP_  (.D(_00249_),
    .DE(_00125_),
    .Q(\w[12][31] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][3]$_DFFE_PP_  (.D(_00250_),
    .DE(_00125_),
    .Q(\w[12][3] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][4]$_DFFE_PP_  (.D(_00251_),
    .DE(_00125_),
    .Q(\w[12][4] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][5]$_DFFE_PP_  (.D(_00252_),
    .DE(_00125_),
    .Q(\w[12][5] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][6]$_DFFE_PP_  (.D(_00253_),
    .DE(_00125_),
    .Q(\w[12][6] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][7]$_DFFE_PP_  (.D(_00254_),
    .DE(_00125_),
    .Q(\w[12][7] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][8]$_DFFE_PP_  (.D(_00255_),
    .DE(_00125_),
    .Q(\w[12][8] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[12][9]$_DFFE_PP_  (.D(_00256_),
    .DE(_00125_),
    .Q(\w[12][9] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][0]$_DFFE_PP_  (.D(_00257_),
    .DE(_00094_),
    .Q(\w[13][0] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][10]$_DFFE_PP_  (.D(_00258_),
    .DE(_00094_),
    .Q(\w[13][10] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][11]$_DFFE_PP_  (.D(_00259_),
    .DE(_00094_),
    .Q(\w[13][11] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][12]$_DFFE_PP_  (.D(_00260_),
    .DE(_00094_),
    .Q(\w[13][12] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][13]$_DFFE_PP_  (.D(_00261_),
    .DE(_00094_),
    .Q(\w[13][13] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][14]$_DFFE_PP_  (.D(_00262_),
    .DE(_00094_),
    .Q(\w[13][14] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][15]$_DFFE_PP_  (.D(_00263_),
    .DE(_00094_),
    .Q(\w[13][15] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][16]$_DFFE_PP_  (.D(_00264_),
    .DE(_00094_),
    .Q(\w[13][16] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][17]$_DFFE_PP_  (.D(_00265_),
    .DE(_00094_),
    .Q(\w[13][17] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][18]$_DFFE_PP_  (.D(_00266_),
    .DE(_00094_),
    .Q(\w[13][18] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][19]$_DFFE_PP_  (.D(_00267_),
    .DE(_00094_),
    .Q(\w[13][19] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][1]$_DFFE_PP_  (.D(_00268_),
    .DE(_00094_),
    .Q(\w[13][1] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][20]$_DFFE_PP_  (.D(_00269_),
    .DE(_00094_),
    .Q(\w[13][20] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][21]$_DFFE_PP_  (.D(_00270_),
    .DE(_00094_),
    .Q(\w[13][21] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][22]$_DFFE_PP_  (.D(_00271_),
    .DE(_00094_),
    .Q(\w[13][22] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][23]$_DFFE_PP_  (.D(_00272_),
    .DE(_00094_),
    .Q(\w[13][23] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][24]$_DFFE_PP_  (.D(_00273_),
    .DE(_00094_),
    .Q(\w[13][24] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][25]$_DFFE_PP_  (.D(_00274_),
    .DE(_00094_),
    .Q(\w[13][25] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][26]$_DFFE_PP_  (.D(_00275_),
    .DE(_00094_),
    .Q(\w[13][26] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][27]$_DFFE_PP_  (.D(_00276_),
    .DE(_00094_),
    .Q(\w[13][27] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][28]$_DFFE_PP_  (.D(_00277_),
    .DE(_00094_),
    .Q(\w[13][28] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][29]$_DFFE_PP_  (.D(_00278_),
    .DE(_00094_),
    .Q(\w[13][29] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][2]$_DFFE_PP_  (.D(_00279_),
    .DE(_00094_),
    .Q(\w[13][2] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][30]$_DFFE_PP_  (.D(_00280_),
    .DE(_00094_),
    .Q(\w[13][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][31]$_DFFE_PP_  (.D(_00281_),
    .DE(_00094_),
    .Q(\w[13][31] ),
    .CLK(clknet_leaf_289_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][3]$_DFFE_PP_  (.D(_00282_),
    .DE(_00094_),
    .Q(\w[13][3] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][4]$_DFFE_PP_  (.D(_00283_),
    .DE(_00094_),
    .Q(\w[13][4] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][5]$_DFFE_PP_  (.D(_00284_),
    .DE(_00094_),
    .Q(\w[13][5] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][6]$_DFFE_PP_  (.D(_00285_),
    .DE(_00094_),
    .Q(\w[13][6] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][7]$_DFFE_PP_  (.D(_00286_),
    .DE(_00094_),
    .Q(\w[13][7] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][8]$_DFFE_PP_  (.D(_00287_),
    .DE(_00094_),
    .Q(\w[13][8] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[13][9]$_DFFE_PP_  (.D(_00288_),
    .DE(_00094_),
    .Q(\w[13][9] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][0]$_DFFE_PP_  (.D(_00289_),
    .DE(_00124_),
    .Q(\w[14][0] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][10]$_DFFE_PP_  (.D(_00290_),
    .DE(_00124_),
    .Q(\w[14][10] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][11]$_DFFE_PP_  (.D(_00291_),
    .DE(_00124_),
    .Q(\w[14][11] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][12]$_DFFE_PP_  (.D(_00292_),
    .DE(_00124_),
    .Q(\w[14][12] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][13]$_DFFE_PP_  (.D(_00293_),
    .DE(_00124_),
    .Q(\w[14][13] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][14]$_DFFE_PP_  (.D(_00294_),
    .DE(_00124_),
    .Q(\w[14][14] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][15]$_DFFE_PP_  (.D(_00295_),
    .DE(_00124_),
    .Q(\w[14][15] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][16]$_DFFE_PP_  (.D(_00296_),
    .DE(_00124_),
    .Q(\w[14][16] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][17]$_DFFE_PP_  (.D(_00297_),
    .DE(_00124_),
    .Q(\w[14][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][18]$_DFFE_PP_  (.D(_00298_),
    .DE(_00124_),
    .Q(\w[14][18] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][19]$_DFFE_PP_  (.D(_00299_),
    .DE(_00124_),
    .Q(\w[14][19] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][1]$_DFFE_PP_  (.D(_00300_),
    .DE(_00124_),
    .Q(\w[14][1] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][20]$_DFFE_PP_  (.D(_00301_),
    .DE(_00124_),
    .Q(\w[14][20] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][21]$_DFFE_PP_  (.D(_00302_),
    .DE(_00124_),
    .Q(\w[14][21] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][22]$_DFFE_PP_  (.D(_00303_),
    .DE(_00124_),
    .Q(\w[14][22] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][23]$_DFFE_PP_  (.D(_00304_),
    .DE(_00124_),
    .Q(\w[14][23] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][24]$_DFFE_PP_  (.D(_00305_),
    .DE(_00124_),
    .Q(\w[14][24] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][25]$_DFFE_PP_  (.D(_00306_),
    .DE(_00124_),
    .Q(\w[14][25] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][26]$_DFFE_PP_  (.D(_00307_),
    .DE(_00124_),
    .Q(\w[14][26] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][27]$_DFFE_PP_  (.D(_00308_),
    .DE(_00124_),
    .Q(\w[14][27] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][28]$_DFFE_PP_  (.D(_00309_),
    .DE(_00124_),
    .Q(\w[14][28] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][29]$_DFFE_PP_  (.D(_00310_),
    .DE(_00124_),
    .Q(\w[14][29] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][2]$_DFFE_PP_  (.D(_00311_),
    .DE(_00124_),
    .Q(\w[14][2] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][30]$_DFFE_PP_  (.D(_00312_),
    .DE(_00124_),
    .Q(\w[14][30] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][31]$_DFFE_PP_  (.D(_00313_),
    .DE(_00124_),
    .Q(\w[14][31] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][3]$_DFFE_PP_  (.D(_00314_),
    .DE(_00124_),
    .Q(\w[14][3] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][4]$_DFFE_PP_  (.D(_00315_),
    .DE(_00124_),
    .Q(\w[14][4] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][5]$_DFFE_PP_  (.D(_00316_),
    .DE(_00124_),
    .Q(\w[14][5] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][6]$_DFFE_PP_  (.D(_00317_),
    .DE(_00124_),
    .Q(\w[14][6] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][7]$_DFFE_PP_  (.D(_00318_),
    .DE(_00124_),
    .Q(\w[14][7] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][8]$_DFFE_PP_  (.D(_00319_),
    .DE(_00124_),
    .Q(\w[14][8] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[14][9]$_DFFE_PP_  (.D(_00320_),
    .DE(_00124_),
    .Q(\w[14][9] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][0]$_DFFE_PP_  (.D(_00321_),
    .DE(_00093_),
    .Q(\w[15][0] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][10]$_DFFE_PP_  (.D(_00322_),
    .DE(_00093_),
    .Q(\w[15][10] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][11]$_DFFE_PP_  (.D(_00323_),
    .DE(_00093_),
    .Q(\w[15][11] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][12]$_DFFE_PP_  (.D(_00324_),
    .DE(_00093_),
    .Q(\w[15][12] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][13]$_DFFE_PP_  (.D(_00325_),
    .DE(_00093_),
    .Q(\w[15][13] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][14]$_DFFE_PP_  (.D(_00326_),
    .DE(_00093_),
    .Q(\w[15][14] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][15]$_DFFE_PP_  (.D(_00327_),
    .DE(_00093_),
    .Q(\w[15][15] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][16]$_DFFE_PP_  (.D(_00328_),
    .DE(_00093_),
    .Q(\w[15][16] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][17]$_DFFE_PP_  (.D(_00329_),
    .DE(_00093_),
    .Q(\w[15][17] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][18]$_DFFE_PP_  (.D(_00330_),
    .DE(_00093_),
    .Q(\w[15][18] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][19]$_DFFE_PP_  (.D(_00331_),
    .DE(_00093_),
    .Q(\w[15][19] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][1]$_DFFE_PP_  (.D(_00332_),
    .DE(_00093_),
    .Q(\w[15][1] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][20]$_DFFE_PP_  (.D(_00333_),
    .DE(_00093_),
    .Q(\w[15][20] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][21]$_DFFE_PP_  (.D(_00334_),
    .DE(_00093_),
    .Q(\w[15][21] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][22]$_DFFE_PP_  (.D(_00335_),
    .DE(_00093_),
    .Q(\w[15][22] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][23]$_DFFE_PP_  (.D(_00336_),
    .DE(_00093_),
    .Q(\w[15][23] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][24]$_DFFE_PP_  (.D(_00337_),
    .DE(_00093_),
    .Q(\w[15][24] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][25]$_DFFE_PP_  (.D(_00338_),
    .DE(_00093_),
    .Q(\w[15][25] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][26]$_DFFE_PP_  (.D(_00339_),
    .DE(_00093_),
    .Q(\w[15][26] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][27]$_DFFE_PP_  (.D(_00340_),
    .DE(_00093_),
    .Q(\w[15][27] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][28]$_DFFE_PP_  (.D(_00341_),
    .DE(_00093_),
    .Q(\w[15][28] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][29]$_DFFE_PP_  (.D(_00342_),
    .DE(_00093_),
    .Q(\w[15][29] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][2]$_DFFE_PP_  (.D(_00343_),
    .DE(_00093_),
    .Q(\w[15][2] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][30]$_DFFE_PP_  (.D(_00344_),
    .DE(_00093_),
    .Q(\w[15][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][31]$_DFFE_PP_  (.D(_00345_),
    .DE(_00093_),
    .Q(\w[15][31] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][3]$_DFFE_PP_  (.D(_00346_),
    .DE(_00093_),
    .Q(\w[15][3] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][4]$_DFFE_PP_  (.D(_00347_),
    .DE(_00093_),
    .Q(\w[15][4] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][5]$_DFFE_PP_  (.D(_00348_),
    .DE(_00093_),
    .Q(\w[15][5] ),
    .CLK(clknet_leaf_290_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][6]$_DFFE_PP_  (.D(_00349_),
    .DE(_00093_),
    .Q(\w[15][6] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][7]$_DFFE_PP_  (.D(_00350_),
    .DE(_00093_),
    .Q(\w[15][7] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][8]$_DFFE_PP_  (.D(_00351_),
    .DE(_00093_),
    .Q(\w[15][8] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[15][9]$_DFFE_PP_  (.D(_00352_),
    .DE(_00093_),
    .Q(\w[15][9] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][0]$_SDFFCE_PN0P_  (.D(_01034_),
    .DE(_00123_),
    .Q(\w[16][0] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][10]$_SDFFCE_PN0P_  (.D(_01035_),
    .DE(_00123_),
    .Q(\w[16][10] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][11]$_SDFFCE_PN0P_  (.D(_01036_),
    .DE(_00123_),
    .Q(\w[16][11] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][12]$_SDFFCE_PN0P_  (.D(_01037_),
    .DE(_00123_),
    .Q(\w[16][12] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][13]$_SDFFCE_PN0P_  (.D(_01038_),
    .DE(_00123_),
    .Q(\w[16][13] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][14]$_SDFFCE_PN0P_  (.D(_01039_),
    .DE(_00123_),
    .Q(\w[16][14] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][15]$_SDFFCE_PN0P_  (.D(_01040_),
    .DE(_00123_),
    .Q(\w[16][15] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][16]$_SDFFCE_PN0P_  (.D(_01041_),
    .DE(_00123_),
    .Q(\w[16][16] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][17]$_SDFFCE_PN0P_  (.D(_01042_),
    .DE(_00123_),
    .Q(\w[16][17] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][18]$_SDFFCE_PN0P_  (.D(_01043_),
    .DE(_00123_),
    .Q(\w[16][18] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][19]$_SDFFCE_PN0P_  (.D(_01044_),
    .DE(_00123_),
    .Q(\w[16][19] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][1]$_SDFFCE_PN0P_  (.D(_01045_),
    .DE(_00123_),
    .Q(\w[16][1] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][20]$_SDFFCE_PN0P_  (.D(_01046_),
    .DE(_00123_),
    .Q(\w[16][20] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][21]$_SDFFCE_PN0P_  (.D(_01047_),
    .DE(_00123_),
    .Q(\w[16][21] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][22]$_SDFFCE_PN0P_  (.D(_01048_),
    .DE(_00123_),
    .Q(\w[16][22] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][23]$_SDFFCE_PN0P_  (.D(_01049_),
    .DE(_00123_),
    .Q(\w[16][23] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][24]$_SDFFCE_PN0P_  (.D(_01050_),
    .DE(_00123_),
    .Q(\w[16][24] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][25]$_SDFFCE_PN0P_  (.D(_01051_),
    .DE(_00123_),
    .Q(\w[16][25] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][26]$_SDFFCE_PN0P_  (.D(_01052_),
    .DE(_00123_),
    .Q(\w[16][26] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][27]$_SDFFCE_PN0P_  (.D(_01053_),
    .DE(_00123_),
    .Q(\w[16][27] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][28]$_SDFFCE_PN0P_  (.D(_01054_),
    .DE(_00123_),
    .Q(\w[16][28] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][29]$_SDFFCE_PN0P_  (.D(_01055_),
    .DE(_00123_),
    .Q(\w[16][29] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][2]$_SDFFCE_PN0P_  (.D(_01056_),
    .DE(_00123_),
    .Q(\w[16][2] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][30]$_SDFFCE_PN0P_  (.D(_01057_),
    .DE(_00123_),
    .Q(\w[16][30] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][31]$_SDFFCE_PN0P_  (.D(_01058_),
    .DE(_00123_),
    .Q(\w[16][31] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][3]$_SDFFCE_PN0P_  (.D(_01059_),
    .DE(_00123_),
    .Q(\w[16][3] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][4]$_SDFFCE_PN0P_  (.D(_01060_),
    .DE(_00123_),
    .Q(\w[16][4] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][5]$_SDFFCE_PN0P_  (.D(_01061_),
    .DE(_00123_),
    .Q(\w[16][5] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][6]$_SDFFCE_PN0P_  (.D(_01062_),
    .DE(_00123_),
    .Q(\w[16][6] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][7]$_SDFFCE_PN0P_  (.D(_01063_),
    .DE(_00123_),
    .Q(\w[16][7] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][8]$_SDFFCE_PN0P_  (.D(_01064_),
    .DE(_00123_),
    .Q(\w[16][8] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[16][9]$_SDFFCE_PN0P_  (.D(_01065_),
    .DE(_00123_),
    .Q(\w[16][9] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][0]$_SDFFCE_PN0P_  (.D(_01066_),
    .DE(_00092_),
    .Q(\w[17][0] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][10]$_SDFFCE_PN0P_  (.D(_01067_),
    .DE(_00092_),
    .Q(\w[17][10] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][11]$_SDFFCE_PN0P_  (.D(_01068_),
    .DE(_00092_),
    .Q(\w[17][11] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][12]$_SDFFCE_PN0P_  (.D(_01069_),
    .DE(_00092_),
    .Q(\w[17][12] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][13]$_SDFFCE_PN0P_  (.D(_01070_),
    .DE(_00092_),
    .Q(\w[17][13] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][14]$_SDFFCE_PN0P_  (.D(_01071_),
    .DE(_00092_),
    .Q(\w[17][14] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][15]$_SDFFCE_PN0P_  (.D(_01072_),
    .DE(_00092_),
    .Q(\w[17][15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][16]$_SDFFCE_PN0P_  (.D(_01073_),
    .DE(_00092_),
    .Q(\w[17][16] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][17]$_SDFFCE_PN0P_  (.D(_01074_),
    .DE(_00092_),
    .Q(\w[17][17] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][18]$_SDFFCE_PN0P_  (.D(_01075_),
    .DE(_00092_),
    .Q(\w[17][18] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][19]$_SDFFCE_PN0P_  (.D(_01076_),
    .DE(_00092_),
    .Q(\w[17][19] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][1]$_SDFFCE_PN0P_  (.D(_01077_),
    .DE(_00092_),
    .Q(\w[17][1] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][20]$_SDFFCE_PN0P_  (.D(_01078_),
    .DE(_00092_),
    .Q(\w[17][20] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][21]$_SDFFCE_PN0P_  (.D(_01079_),
    .DE(_00092_),
    .Q(\w[17][21] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][22]$_SDFFCE_PN0P_  (.D(_01080_),
    .DE(_00092_),
    .Q(\w[17][22] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][23]$_SDFFCE_PN0P_  (.D(_01081_),
    .DE(_00092_),
    .Q(\w[17][23] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][24]$_SDFFCE_PN0P_  (.D(_01082_),
    .DE(_00092_),
    .Q(\w[17][24] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][25]$_SDFFCE_PN0P_  (.D(_01083_),
    .DE(_00092_),
    .Q(\w[17][25] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][26]$_SDFFCE_PN0P_  (.D(_01084_),
    .DE(_00092_),
    .Q(\w[17][26] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][27]$_SDFFCE_PN0P_  (.D(_01085_),
    .DE(_00092_),
    .Q(\w[17][27] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][28]$_SDFFCE_PN0P_  (.D(_01086_),
    .DE(_00092_),
    .Q(\w[17][28] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][29]$_SDFFCE_PN0P_  (.D(_01087_),
    .DE(_00092_),
    .Q(\w[17][29] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][2]$_SDFFCE_PN0P_  (.D(_01088_),
    .DE(_00092_),
    .Q(\w[17][2] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][30]$_SDFFCE_PN0P_  (.D(_01089_),
    .DE(_00092_),
    .Q(\w[17][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][31]$_SDFFCE_PN0P_  (.D(_01090_),
    .DE(_00092_),
    .Q(\w[17][31] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][3]$_SDFFCE_PN0P_  (.D(_01091_),
    .DE(_00092_),
    .Q(\w[17][3] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][4]$_SDFFCE_PN0P_  (.D(_01092_),
    .DE(_00092_),
    .Q(\w[17][4] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][5]$_SDFFCE_PN0P_  (.D(_01093_),
    .DE(_00092_),
    .Q(\w[17][5] ),
    .CLK(clknet_leaf_290_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][6]$_SDFFCE_PN0P_  (.D(_01094_),
    .DE(_00092_),
    .Q(\w[17][6] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][7]$_SDFFCE_PN0P_  (.D(_01095_),
    .DE(_00092_),
    .Q(\w[17][7] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][8]$_SDFFCE_PN0P_  (.D(_01096_),
    .DE(_00092_),
    .Q(\w[17][8] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[17][9]$_SDFFCE_PN0P_  (.D(_01097_),
    .DE(_00092_),
    .Q(\w[17][9] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][0]$_SDFFCE_PN0P_  (.D(_01098_),
    .DE(_00122_),
    .Q(\w[18][0] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][10]$_SDFFCE_PN0P_  (.D(_01099_),
    .DE(_00122_),
    .Q(\w[18][10] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][11]$_SDFFCE_PN0P_  (.D(_01100_),
    .DE(_00122_),
    .Q(\w[18][11] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][12]$_SDFFCE_PN0P_  (.D(_01101_),
    .DE(_00122_),
    .Q(\w[18][12] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][13]$_SDFFCE_PN0P_  (.D(_01102_),
    .DE(_00122_),
    .Q(\w[18][13] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][14]$_SDFFCE_PN0P_  (.D(_01103_),
    .DE(_00122_),
    .Q(\w[18][14] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][15]$_SDFFCE_PN0P_  (.D(_01104_),
    .DE(_00122_),
    .Q(\w[18][15] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][16]$_SDFFCE_PN0P_  (.D(_01105_),
    .DE(_00122_),
    .Q(\w[18][16] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][17]$_SDFFCE_PN0P_  (.D(_01106_),
    .DE(_00122_),
    .Q(\w[18][17] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][18]$_SDFFCE_PN0P_  (.D(_01107_),
    .DE(_00122_),
    .Q(\w[18][18] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][19]$_SDFFCE_PN0P_  (.D(_01108_),
    .DE(_00122_),
    .Q(\w[18][19] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][1]$_SDFFCE_PN0P_  (.D(_01109_),
    .DE(_00122_),
    .Q(\w[18][1] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][20]$_SDFFCE_PN0P_  (.D(_01110_),
    .DE(_00122_),
    .Q(\w[18][20] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][21]$_SDFFCE_PN0P_  (.D(_01111_),
    .DE(_00122_),
    .Q(\w[18][21] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][22]$_SDFFCE_PN0P_  (.D(_01112_),
    .DE(_00122_),
    .Q(\w[18][22] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][23]$_SDFFCE_PN0P_  (.D(_01113_),
    .DE(_00122_),
    .Q(\w[18][23] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][24]$_SDFFCE_PN0P_  (.D(_01114_),
    .DE(_00122_),
    .Q(\w[18][24] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][25]$_SDFFCE_PN0P_  (.D(_01115_),
    .DE(_00122_),
    .Q(\w[18][25] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][26]$_SDFFCE_PN0P_  (.D(_01116_),
    .DE(_00122_),
    .Q(\w[18][26] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][27]$_SDFFCE_PN0P_  (.D(_01117_),
    .DE(_00122_),
    .Q(\w[18][27] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][28]$_SDFFCE_PN0P_  (.D(_01118_),
    .DE(_00122_),
    .Q(\w[18][28] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][29]$_SDFFCE_PN0P_  (.D(_01119_),
    .DE(_00122_),
    .Q(\w[18][29] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][2]$_SDFFCE_PN0P_  (.D(_01120_),
    .DE(_00122_),
    .Q(\w[18][2] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][30]$_SDFFCE_PN0P_  (.D(_01121_),
    .DE(_00122_),
    .Q(\w[18][30] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][31]$_SDFFCE_PN0P_  (.D(_01122_),
    .DE(_00122_),
    .Q(\w[18][31] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][3]$_SDFFCE_PN0P_  (.D(_01123_),
    .DE(_00122_),
    .Q(\w[18][3] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][4]$_SDFFCE_PN0P_  (.D(_01124_),
    .DE(_00122_),
    .Q(\w[18][4] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][5]$_SDFFCE_PN0P_  (.D(_01125_),
    .DE(_00122_),
    .Q(\w[18][5] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][6]$_SDFFCE_PN0P_  (.D(_01126_),
    .DE(_00122_),
    .Q(\w[18][6] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][7]$_SDFFCE_PN0P_  (.D(_01127_),
    .DE(_00122_),
    .Q(\w[18][7] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][8]$_SDFFCE_PN0P_  (.D(_01128_),
    .DE(_00122_),
    .Q(\w[18][8] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[18][9]$_SDFFCE_PN0P_  (.D(_01129_),
    .DE(_00122_),
    .Q(\w[18][9] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][0]$_SDFFCE_PN0P_  (.D(_01130_),
    .DE(_00091_),
    .Q(\w[19][0] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][10]$_SDFFCE_PN0P_  (.D(_01131_),
    .DE(_00091_),
    .Q(\w[19][10] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][11]$_SDFFCE_PN0P_  (.D(_01132_),
    .DE(_00091_),
    .Q(\w[19][11] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][12]$_SDFFCE_PN0P_  (.D(_01133_),
    .DE(_00091_),
    .Q(\w[19][12] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][13]$_SDFFCE_PN0P_  (.D(_01134_),
    .DE(_00091_),
    .Q(\w[19][13] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][14]$_SDFFCE_PN0P_  (.D(_01135_),
    .DE(_00091_),
    .Q(\w[19][14] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][15]$_SDFFCE_PN0P_  (.D(_01136_),
    .DE(_00091_),
    .Q(\w[19][15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][16]$_SDFFCE_PN0P_  (.D(_01137_),
    .DE(_00091_),
    .Q(\w[19][16] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][17]$_SDFFCE_PN0P_  (.D(_01138_),
    .DE(_00091_),
    .Q(\w[19][17] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][18]$_SDFFCE_PN0P_  (.D(_01139_),
    .DE(_00091_),
    .Q(\w[19][18] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][19]$_SDFFCE_PN0P_  (.D(_01140_),
    .DE(_00091_),
    .Q(\w[19][19] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][1]$_SDFFCE_PN0P_  (.D(_01141_),
    .DE(_00091_),
    .Q(\w[19][1] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][20]$_SDFFCE_PN0P_  (.D(_01142_),
    .DE(_00091_),
    .Q(\w[19][20] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][21]$_SDFFCE_PN0P_  (.D(_01143_),
    .DE(_00091_),
    .Q(\w[19][21] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][22]$_SDFFCE_PN0P_  (.D(_01144_),
    .DE(_00091_),
    .Q(\w[19][22] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][23]$_SDFFCE_PN0P_  (.D(_01145_),
    .DE(_00091_),
    .Q(\w[19][23] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][24]$_SDFFCE_PN0P_  (.D(_01146_),
    .DE(_00091_),
    .Q(\w[19][24] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][25]$_SDFFCE_PN0P_  (.D(_01147_),
    .DE(_00091_),
    .Q(\w[19][25] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][26]$_SDFFCE_PN0P_  (.D(_01148_),
    .DE(_00091_),
    .Q(\w[19][26] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][27]$_SDFFCE_PN0P_  (.D(_01149_),
    .DE(_00091_),
    .Q(\w[19][27] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][28]$_SDFFCE_PN0P_  (.D(_01150_),
    .DE(_00091_),
    .Q(\w[19][28] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][29]$_SDFFCE_PN0P_  (.D(_01151_),
    .DE(_00091_),
    .Q(\w[19][29] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][2]$_SDFFCE_PN0P_  (.D(_01152_),
    .DE(_00091_),
    .Q(\w[19][2] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][30]$_SDFFCE_PN0P_  (.D(_01153_),
    .DE(_00091_),
    .Q(\w[19][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][31]$_SDFFCE_PN0P_  (.D(_01154_),
    .DE(_00091_),
    .Q(\w[19][31] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][3]$_SDFFCE_PN0P_  (.D(_01155_),
    .DE(_00091_),
    .Q(\w[19][3] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][4]$_SDFFCE_PN0P_  (.D(_01156_),
    .DE(_00091_),
    .Q(\w[19][4] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][5]$_SDFFCE_PN0P_  (.D(_01157_),
    .DE(_00091_),
    .Q(\w[19][5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][6]$_SDFFCE_PN0P_  (.D(_01158_),
    .DE(_00091_),
    .Q(\w[19][6] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][7]$_SDFFCE_PN0P_  (.D(_01159_),
    .DE(_00091_),
    .Q(\w[19][7] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][8]$_SDFFCE_PN0P_  (.D(_01160_),
    .DE(_00091_),
    .Q(\w[19][8] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[19][9]$_SDFFCE_PN0P_  (.D(_01161_),
    .DE(_00091_),
    .Q(\w[19][9] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][0]$_DFFE_PP_  (.D(_00353_),
    .DE(_00090_),
    .Q(\w[1][0] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][10]$_DFFE_PP_  (.D(_00354_),
    .DE(_00090_),
    .Q(\w[1][10] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][11]$_DFFE_PP_  (.D(_00355_),
    .DE(_00090_),
    .Q(\w[1][11] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][12]$_DFFE_PP_  (.D(_00356_),
    .DE(_00090_),
    .Q(\w[1][12] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][13]$_DFFE_PP_  (.D(_00357_),
    .DE(_00090_),
    .Q(\w[1][13] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][14]$_DFFE_PP_  (.D(_00358_),
    .DE(_00090_),
    .Q(\w[1][14] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][15]$_DFFE_PP_  (.D(_00359_),
    .DE(_00090_),
    .Q(\w[1][15] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][16]$_DFFE_PP_  (.D(_00360_),
    .DE(_00090_),
    .Q(\w[1][16] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][17]$_DFFE_PP_  (.D(_00361_),
    .DE(_00090_),
    .Q(\w[1][17] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][18]$_DFFE_PP_  (.D(_00362_),
    .DE(_00090_),
    .Q(\w[1][18] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][19]$_DFFE_PP_  (.D(_00363_),
    .DE(_00090_),
    .Q(\w[1][19] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][1]$_DFFE_PP_  (.D(_00364_),
    .DE(_00090_),
    .Q(\w[1][1] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][20]$_DFFE_PP_  (.D(_00365_),
    .DE(_00090_),
    .Q(\w[1][20] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][21]$_DFFE_PP_  (.D(_00366_),
    .DE(_00090_),
    .Q(\w[1][21] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][22]$_DFFE_PP_  (.D(_00367_),
    .DE(_00090_),
    .Q(\w[1][22] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][23]$_DFFE_PP_  (.D(_00368_),
    .DE(_00090_),
    .Q(\w[1][23] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][24]$_DFFE_PP_  (.D(_00369_),
    .DE(_00090_),
    .Q(\w[1][24] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][25]$_DFFE_PP_  (.D(_00370_),
    .DE(_00090_),
    .Q(\w[1][25] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][26]$_DFFE_PP_  (.D(_00371_),
    .DE(_00090_),
    .Q(\w[1][26] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][27]$_DFFE_PP_  (.D(_00372_),
    .DE(_00090_),
    .Q(\w[1][27] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][28]$_DFFE_PP_  (.D(_00373_),
    .DE(_00090_),
    .Q(\w[1][28] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][29]$_DFFE_PP_  (.D(_00374_),
    .DE(_00090_),
    .Q(\w[1][29] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][2]$_DFFE_PP_  (.D(_00375_),
    .DE(_00090_),
    .Q(\w[1][2] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][30]$_DFFE_PP_  (.D(_00376_),
    .DE(_00090_),
    .Q(\w[1][30] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][31]$_DFFE_PP_  (.D(_00377_),
    .DE(_00090_),
    .Q(\w[1][31] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][3]$_DFFE_PP_  (.D(_00378_),
    .DE(_00090_),
    .Q(\w[1][3] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][4]$_DFFE_PP_  (.D(_00379_),
    .DE(_00090_),
    .Q(\w[1][4] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][5]$_DFFE_PP_  (.D(_00380_),
    .DE(_00090_),
    .Q(\w[1][5] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][6]$_DFFE_PP_  (.D(_00381_),
    .DE(_00090_),
    .Q(\w[1][6] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][7]$_DFFE_PP_  (.D(_00382_),
    .DE(_00090_),
    .Q(\w[1][7] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][8]$_DFFE_PP_  (.D(_00383_),
    .DE(_00090_),
    .Q(\w[1][8] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[1][9]$_DFFE_PP_  (.D(_00384_),
    .DE(_00090_),
    .Q(\w[1][9] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][0]$_SDFFCE_PN0P_  (.D(_01162_),
    .DE(_00121_),
    .Q(\w[20][0] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][10]$_SDFFCE_PN0P_  (.D(_01163_),
    .DE(_00121_),
    .Q(\w[20][10] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][11]$_SDFFCE_PN0P_  (.D(_01164_),
    .DE(_00121_),
    .Q(\w[20][11] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][12]$_SDFFCE_PN0P_  (.D(_01165_),
    .DE(_00121_),
    .Q(\w[20][12] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][13]$_SDFFCE_PN0P_  (.D(_01166_),
    .DE(_00121_),
    .Q(\w[20][13] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][14]$_SDFFCE_PN0P_  (.D(_01167_),
    .DE(_00121_),
    .Q(\w[20][14] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][15]$_SDFFCE_PN0P_  (.D(_01168_),
    .DE(_00121_),
    .Q(\w[20][15] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][16]$_SDFFCE_PN0P_  (.D(_01169_),
    .DE(_00121_),
    .Q(\w[20][16] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][17]$_SDFFCE_PN0P_  (.D(_01170_),
    .DE(_00121_),
    .Q(\w[20][17] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][18]$_SDFFCE_PN0P_  (.D(_01171_),
    .DE(_00121_),
    .Q(\w[20][18] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][19]$_SDFFCE_PN0P_  (.D(_01172_),
    .DE(_00121_),
    .Q(\w[20][19] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][1]$_SDFFCE_PN0P_  (.D(_01173_),
    .DE(_00121_),
    .Q(\w[20][1] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][20]$_SDFFCE_PN0P_  (.D(_01174_),
    .DE(_00121_),
    .Q(\w[20][20] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][21]$_SDFFCE_PN0P_  (.D(_01175_),
    .DE(_00121_),
    .Q(\w[20][21] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][22]$_SDFFCE_PN0P_  (.D(_01176_),
    .DE(_00121_),
    .Q(\w[20][22] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][23]$_SDFFCE_PN0P_  (.D(_01177_),
    .DE(_00121_),
    .Q(\w[20][23] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][24]$_SDFFCE_PN0P_  (.D(_01178_),
    .DE(_00121_),
    .Q(\w[20][24] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][25]$_SDFFCE_PN0P_  (.D(_01179_),
    .DE(_00121_),
    .Q(\w[20][25] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][26]$_SDFFCE_PN0P_  (.D(_01180_),
    .DE(_00121_),
    .Q(\w[20][26] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][27]$_SDFFCE_PN0P_  (.D(_01181_),
    .DE(_00121_),
    .Q(\w[20][27] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][28]$_SDFFCE_PN0P_  (.D(_01182_),
    .DE(_00121_),
    .Q(\w[20][28] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][29]$_SDFFCE_PN0P_  (.D(_01183_),
    .DE(_00121_),
    .Q(\w[20][29] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][2]$_SDFFCE_PN0P_  (.D(_01184_),
    .DE(_00121_),
    .Q(\w[20][2] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][30]$_SDFFCE_PN0P_  (.D(_01185_),
    .DE(_00121_),
    .Q(\w[20][30] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][31]$_SDFFCE_PN0P_  (.D(_01186_),
    .DE(_00121_),
    .Q(\w[20][31] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][3]$_SDFFCE_PN0P_  (.D(_01187_),
    .DE(_00121_),
    .Q(\w[20][3] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][4]$_SDFFCE_PN0P_  (.D(_01188_),
    .DE(_00121_),
    .Q(\w[20][4] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][5]$_SDFFCE_PN0P_  (.D(_01189_),
    .DE(_00121_),
    .Q(\w[20][5] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][6]$_SDFFCE_PN0P_  (.D(_01190_),
    .DE(_00121_),
    .Q(\w[20][6] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][7]$_SDFFCE_PN0P_  (.D(_01191_),
    .DE(_00121_),
    .Q(\w[20][7] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][8]$_SDFFCE_PN0P_  (.D(_01192_),
    .DE(_00121_),
    .Q(\w[20][8] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[20][9]$_SDFFCE_PN0P_  (.D(_01193_),
    .DE(_00121_),
    .Q(\w[20][9] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][0]$_SDFFCE_PN0P_  (.D(_01194_),
    .DE(_00089_),
    .Q(\w[21][0] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][10]$_SDFFCE_PN0P_  (.D(_01195_),
    .DE(_00089_),
    .Q(\w[21][10] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][11]$_SDFFCE_PN0P_  (.D(_01196_),
    .DE(_00089_),
    .Q(\w[21][11] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][12]$_SDFFCE_PN0P_  (.D(_01197_),
    .DE(_00089_),
    .Q(\w[21][12] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][13]$_SDFFCE_PN0P_  (.D(_01198_),
    .DE(_00089_),
    .Q(\w[21][13] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][14]$_SDFFCE_PN0P_  (.D(_01199_),
    .DE(_00089_),
    .Q(\w[21][14] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][15]$_SDFFCE_PN0P_  (.D(_01200_),
    .DE(_00089_),
    .Q(\w[21][15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][16]$_SDFFCE_PN0P_  (.D(_01201_),
    .DE(_00089_),
    .Q(\w[21][16] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][17]$_SDFFCE_PN0P_  (.D(_01202_),
    .DE(_00089_),
    .Q(\w[21][17] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][18]$_SDFFCE_PN0P_  (.D(_01203_),
    .DE(_00089_),
    .Q(\w[21][18] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][19]$_SDFFCE_PN0P_  (.D(_01204_),
    .DE(_00089_),
    .Q(\w[21][19] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][1]$_SDFFCE_PN0P_  (.D(_01205_),
    .DE(_00089_),
    .Q(\w[21][1] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][20]$_SDFFCE_PN0P_  (.D(_01206_),
    .DE(_00089_),
    .Q(\w[21][20] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][21]$_SDFFCE_PN0P_  (.D(_01207_),
    .DE(_00089_),
    .Q(\w[21][21] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][22]$_SDFFCE_PN0P_  (.D(_01208_),
    .DE(_00089_),
    .Q(\w[21][22] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][23]$_SDFFCE_PN0P_  (.D(_01209_),
    .DE(_00089_),
    .Q(\w[21][23] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][24]$_SDFFCE_PN0P_  (.D(_01210_),
    .DE(_00089_),
    .Q(\w[21][24] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][25]$_SDFFCE_PN0P_  (.D(_01211_),
    .DE(_00089_),
    .Q(\w[21][25] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][26]$_SDFFCE_PN0P_  (.D(_01212_),
    .DE(_00089_),
    .Q(\w[21][26] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][27]$_SDFFCE_PN0P_  (.D(_01213_),
    .DE(_00089_),
    .Q(\w[21][27] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][28]$_SDFFCE_PN0P_  (.D(_01214_),
    .DE(_00089_),
    .Q(\w[21][28] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][29]$_SDFFCE_PN0P_  (.D(_01215_),
    .DE(_00089_),
    .Q(\w[21][29] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][2]$_SDFFCE_PN0P_  (.D(_01216_),
    .DE(_00089_),
    .Q(\w[21][2] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][30]$_SDFFCE_PN0P_  (.D(_01217_),
    .DE(_00089_),
    .Q(\w[21][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][31]$_SDFFCE_PN0P_  (.D(_01218_),
    .DE(_00089_),
    .Q(\w[21][31] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][3]$_SDFFCE_PN0P_  (.D(_01219_),
    .DE(_00089_),
    .Q(\w[21][3] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][4]$_SDFFCE_PN0P_  (.D(_01220_),
    .DE(_00089_),
    .Q(\w[21][4] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][5]$_SDFFCE_PN0P_  (.D(_01221_),
    .DE(_00089_),
    .Q(\w[21][5] ),
    .CLK(clknet_leaf_290_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][6]$_SDFFCE_PN0P_  (.D(_01222_),
    .DE(_00089_),
    .Q(\w[21][6] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][7]$_SDFFCE_PN0P_  (.D(_01223_),
    .DE(_00089_),
    .Q(\w[21][7] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][8]$_SDFFCE_PN0P_  (.D(_01224_),
    .DE(_00089_),
    .Q(\w[21][8] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[21][9]$_SDFFCE_PN0P_  (.D(_01225_),
    .DE(_00089_),
    .Q(\w[21][9] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][0]$_SDFFCE_PN0P_  (.D(_01226_),
    .DE(_00120_),
    .Q(\w[22][0] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][10]$_SDFFCE_PN0P_  (.D(_01227_),
    .DE(_00120_),
    .Q(\w[22][10] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][11]$_SDFFCE_PN0P_  (.D(_01228_),
    .DE(_00120_),
    .Q(\w[22][11] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][12]$_SDFFCE_PN0P_  (.D(_01229_),
    .DE(_00120_),
    .Q(\w[22][12] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][13]$_SDFFCE_PN0P_  (.D(_01230_),
    .DE(_00120_),
    .Q(\w[22][13] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][14]$_SDFFCE_PN0P_  (.D(_01231_),
    .DE(_00120_),
    .Q(\w[22][14] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][15]$_SDFFCE_PN0P_  (.D(_01232_),
    .DE(_00120_),
    .Q(\w[22][15] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][16]$_SDFFCE_PN0P_  (.D(_01233_),
    .DE(_00120_),
    .Q(\w[22][16] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][17]$_SDFFCE_PN0P_  (.D(_01234_),
    .DE(_00120_),
    .Q(\w[22][17] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][18]$_SDFFCE_PN0P_  (.D(_01235_),
    .DE(_00120_),
    .Q(\w[22][18] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][19]$_SDFFCE_PN0P_  (.D(_01236_),
    .DE(_00120_),
    .Q(\w[22][19] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][1]$_SDFFCE_PN0P_  (.D(_01237_),
    .DE(_00120_),
    .Q(\w[22][1] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][20]$_SDFFCE_PN0P_  (.D(_01238_),
    .DE(_00120_),
    .Q(\w[22][20] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][21]$_SDFFCE_PN0P_  (.D(_01239_),
    .DE(_00120_),
    .Q(\w[22][21] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][22]$_SDFFCE_PN0P_  (.D(_01240_),
    .DE(_00120_),
    .Q(\w[22][22] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][23]$_SDFFCE_PN0P_  (.D(_01241_),
    .DE(_00120_),
    .Q(\w[22][23] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][24]$_SDFFCE_PN0P_  (.D(_01242_),
    .DE(_00120_),
    .Q(\w[22][24] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][25]$_SDFFCE_PN0P_  (.D(_01243_),
    .DE(_00120_),
    .Q(\w[22][25] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][26]$_SDFFCE_PN0P_  (.D(_01244_),
    .DE(_00120_),
    .Q(\w[22][26] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][27]$_SDFFCE_PN0P_  (.D(_01245_),
    .DE(_00120_),
    .Q(\w[22][27] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][28]$_SDFFCE_PN0P_  (.D(_01246_),
    .DE(_00120_),
    .Q(\w[22][28] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][29]$_SDFFCE_PN0P_  (.D(_01247_),
    .DE(_00120_),
    .Q(\w[22][29] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][2]$_SDFFCE_PN0P_  (.D(_01248_),
    .DE(_00120_),
    .Q(\w[22][2] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][30]$_SDFFCE_PN0P_  (.D(_01249_),
    .DE(_00120_),
    .Q(\w[22][30] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][31]$_SDFFCE_PN0P_  (.D(_01250_),
    .DE(_00120_),
    .Q(\w[22][31] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][3]$_SDFFCE_PN0P_  (.D(_01251_),
    .DE(_00120_),
    .Q(\w[22][3] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][4]$_SDFFCE_PN0P_  (.D(_01252_),
    .DE(_00120_),
    .Q(\w[22][4] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][5]$_SDFFCE_PN0P_  (.D(_01253_),
    .DE(_00120_),
    .Q(\w[22][5] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][6]$_SDFFCE_PN0P_  (.D(_01254_),
    .DE(_00120_),
    .Q(\w[22][6] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][7]$_SDFFCE_PN0P_  (.D(_01255_),
    .DE(_00120_),
    .Q(\w[22][7] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][8]$_SDFFCE_PN0P_  (.D(_01256_),
    .DE(_00120_),
    .Q(\w[22][8] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[22][9]$_SDFFCE_PN0P_  (.D(_01257_),
    .DE(_00120_),
    .Q(\w[22][9] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][0]$_SDFFCE_PN0P_  (.D(_01258_),
    .DE(net301),
    .Q(\w[23][0] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][10]$_SDFFCE_PN0P_  (.D(_01259_),
    .DE(net301),
    .Q(\w[23][10] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][11]$_SDFFCE_PN0P_  (.D(_01260_),
    .DE(net301),
    .Q(\w[23][11] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][12]$_SDFFCE_PN0P_  (.D(_01261_),
    .DE(net301),
    .Q(\w[23][12] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][13]$_SDFFCE_PN0P_  (.D(_01262_),
    .DE(net301),
    .Q(\w[23][13] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][14]$_SDFFCE_PN0P_  (.D(_01263_),
    .DE(net301),
    .Q(\w[23][14] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][15]$_SDFFCE_PN0P_  (.D(_01264_),
    .DE(_00088_),
    .Q(\w[23][15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][16]$_SDFFCE_PN0P_  (.D(_01265_),
    .DE(net302),
    .Q(\w[23][16] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][17]$_SDFFCE_PN0P_  (.D(_01266_),
    .DE(net301),
    .Q(\w[23][17] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][18]$_SDFFCE_PN0P_  (.D(_01267_),
    .DE(net301),
    .Q(\w[23][18] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][19]$_SDFFCE_PN0P_  (.D(_01268_),
    .DE(net301),
    .Q(\w[23][19] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][1]$_SDFFCE_PN0P_  (.D(_01269_),
    .DE(net302),
    .Q(\w[23][1] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][20]$_SDFFCE_PN0P_  (.D(_01270_),
    .DE(net301),
    .Q(\w[23][20] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][21]$_SDFFCE_PN0P_  (.D(_01271_),
    .DE(net301),
    .Q(\w[23][21] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][22]$_SDFFCE_PN0P_  (.D(_01272_),
    .DE(net301),
    .Q(\w[23][22] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][23]$_SDFFCE_PN0P_  (.D(_01273_),
    .DE(net302),
    .Q(\w[23][23] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][24]$_SDFFCE_PN0P_  (.D(_01274_),
    .DE(net302),
    .Q(\w[23][24] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][25]$_SDFFCE_PN0P_  (.D(_01275_),
    .DE(net301),
    .Q(\w[23][25] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][26]$_SDFFCE_PN0P_  (.D(_01276_),
    .DE(net302),
    .Q(\w[23][26] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][27]$_SDFFCE_PN0P_  (.D(_01277_),
    .DE(net302),
    .Q(\w[23][27] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][28]$_SDFFCE_PN0P_  (.D(_01278_),
    .DE(net302),
    .Q(\w[23][28] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][29]$_SDFFCE_PN0P_  (.D(_01279_),
    .DE(_00088_),
    .Q(\w[23][29] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][2]$_SDFFCE_PN0P_  (.D(_01280_),
    .DE(net301),
    .Q(\w[23][2] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][30]$_SDFFCE_PN0P_  (.D(_01281_),
    .DE(_00088_),
    .Q(\w[23][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][31]$_SDFFCE_PN0P_  (.D(_01282_),
    .DE(net302),
    .Q(\w[23][31] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][3]$_SDFFCE_PN0P_  (.D(_01283_),
    .DE(net302),
    .Q(\w[23][3] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][4]$_SDFFCE_PN0P_  (.D(_01284_),
    .DE(net302),
    .Q(\w[23][4] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][5]$_SDFFCE_PN0P_  (.D(_01285_),
    .DE(net302),
    .Q(\w[23][5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][6]$_SDFFCE_PN0P_  (.D(_01286_),
    .DE(net302),
    .Q(\w[23][6] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][7]$_SDFFCE_PN0P_  (.D(_01287_),
    .DE(net302),
    .Q(\w[23][7] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][8]$_SDFFCE_PN0P_  (.D(_01288_),
    .DE(net301),
    .Q(\w[23][8] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[23][9]$_SDFFCE_PN0P_  (.D(_01289_),
    .DE(_00088_),
    .Q(\w[23][9] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][0]$_SDFFCE_PN0P_  (.D(_01290_),
    .DE(_00119_),
    .Q(\w[24][0] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][10]$_SDFFCE_PN0P_  (.D(_01291_),
    .DE(_00119_),
    .Q(\w[24][10] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][11]$_SDFFCE_PN0P_  (.D(_01292_),
    .DE(_00119_),
    .Q(\w[24][11] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][12]$_SDFFCE_PN0P_  (.D(_01293_),
    .DE(_00119_),
    .Q(\w[24][12] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][13]$_SDFFCE_PN0P_  (.D(_01294_),
    .DE(_00119_),
    .Q(\w[24][13] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][14]$_SDFFCE_PN0P_  (.D(_01295_),
    .DE(_00119_),
    .Q(\w[24][14] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][15]$_SDFFCE_PN0P_  (.D(_01296_),
    .DE(_00119_),
    .Q(\w[24][15] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][16]$_SDFFCE_PN0P_  (.D(_01297_),
    .DE(_00119_),
    .Q(\w[24][16] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][17]$_SDFFCE_PN0P_  (.D(_01298_),
    .DE(_00119_),
    .Q(\w[24][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][18]$_SDFFCE_PN0P_  (.D(_01299_),
    .DE(_00119_),
    .Q(\w[24][18] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][19]$_SDFFCE_PN0P_  (.D(_01300_),
    .DE(_00119_),
    .Q(\w[24][19] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][1]$_SDFFCE_PN0P_  (.D(_01301_),
    .DE(_00119_),
    .Q(\w[24][1] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][20]$_SDFFCE_PN0P_  (.D(_01302_),
    .DE(_00119_),
    .Q(\w[24][20] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][21]$_SDFFCE_PN0P_  (.D(_01303_),
    .DE(_00119_),
    .Q(\w[24][21] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][22]$_SDFFCE_PN0P_  (.D(_01304_),
    .DE(_00119_),
    .Q(\w[24][22] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][23]$_SDFFCE_PN0P_  (.D(_01305_),
    .DE(_00119_),
    .Q(\w[24][23] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][24]$_SDFFCE_PN0P_  (.D(_01306_),
    .DE(_00119_),
    .Q(\w[24][24] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][25]$_SDFFCE_PN0P_  (.D(_01307_),
    .DE(_00119_),
    .Q(\w[24][25] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][26]$_SDFFCE_PN0P_  (.D(_01308_),
    .DE(_00119_),
    .Q(\w[24][26] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][27]$_SDFFCE_PN0P_  (.D(_01309_),
    .DE(_00119_),
    .Q(\w[24][27] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][28]$_SDFFCE_PN0P_  (.D(_01310_),
    .DE(_00119_),
    .Q(\w[24][28] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][29]$_SDFFCE_PN0P_  (.D(_01311_),
    .DE(_00119_),
    .Q(\w[24][29] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][2]$_SDFFCE_PN0P_  (.D(_01312_),
    .DE(_00119_),
    .Q(\w[24][2] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][30]$_SDFFCE_PN0P_  (.D(_01313_),
    .DE(_00119_),
    .Q(\w[24][30] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][31]$_SDFFCE_PN0P_  (.D(_01314_),
    .DE(_00119_),
    .Q(\w[24][31] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][3]$_SDFFCE_PN0P_  (.D(_01315_),
    .DE(_00119_),
    .Q(\w[24][3] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][4]$_SDFFCE_PN0P_  (.D(_01316_),
    .DE(_00119_),
    .Q(\w[24][4] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][5]$_SDFFCE_PN0P_  (.D(_01317_),
    .DE(_00119_),
    .Q(\w[24][5] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][6]$_SDFFCE_PN0P_  (.D(_01318_),
    .DE(_00119_),
    .Q(\w[24][6] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][7]$_SDFFCE_PN0P_  (.D(_01319_),
    .DE(_00119_),
    .Q(\w[24][7] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][8]$_SDFFCE_PN0P_  (.D(_01320_),
    .DE(_00119_),
    .Q(\w[24][8] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[24][9]$_SDFFCE_PN0P_  (.D(_01321_),
    .DE(_00119_),
    .Q(\w[24][9] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][0]$_SDFFCE_PN0P_  (.D(_01322_),
    .DE(_00087_),
    .Q(\w[25][0] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][10]$_SDFFCE_PN0P_  (.D(_01323_),
    .DE(_00087_),
    .Q(\w[25][10] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][11]$_SDFFCE_PN0P_  (.D(_01324_),
    .DE(_00087_),
    .Q(\w[25][11] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][12]$_SDFFCE_PN0P_  (.D(_01325_),
    .DE(_00087_),
    .Q(\w[25][12] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][13]$_SDFFCE_PN0P_  (.D(_01326_),
    .DE(_00087_),
    .Q(\w[25][13] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][14]$_SDFFCE_PN0P_  (.D(_01327_),
    .DE(_00087_),
    .Q(\w[25][14] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][15]$_SDFFCE_PN0P_  (.D(_01328_),
    .DE(_00087_),
    .Q(\w[25][15] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][16]$_SDFFCE_PN0P_  (.D(_01329_),
    .DE(_00087_),
    .Q(\w[25][16] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][17]$_SDFFCE_PN0P_  (.D(_01330_),
    .DE(_00087_),
    .Q(\w[25][17] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][18]$_SDFFCE_PN0P_  (.D(_01331_),
    .DE(_00087_),
    .Q(\w[25][18] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][19]$_SDFFCE_PN0P_  (.D(_01332_),
    .DE(_00087_),
    .Q(\w[25][19] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][1]$_SDFFCE_PN0P_  (.D(_01333_),
    .DE(_00087_),
    .Q(\w[25][1] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][20]$_SDFFCE_PN0P_  (.D(_01334_),
    .DE(_00087_),
    .Q(\w[25][20] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][21]$_SDFFCE_PN0P_  (.D(_01335_),
    .DE(_00087_),
    .Q(\w[25][21] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][22]$_SDFFCE_PN0P_  (.D(_01336_),
    .DE(_00087_),
    .Q(\w[25][22] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][23]$_SDFFCE_PN0P_  (.D(_01337_),
    .DE(_00087_),
    .Q(\w[25][23] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][24]$_SDFFCE_PN0P_  (.D(_01338_),
    .DE(_00087_),
    .Q(\w[25][24] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][25]$_SDFFCE_PN0P_  (.D(_01339_),
    .DE(_00087_),
    .Q(\w[25][25] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][26]$_SDFFCE_PN0P_  (.D(_01340_),
    .DE(_00087_),
    .Q(\w[25][26] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][27]$_SDFFCE_PN0P_  (.D(_01341_),
    .DE(_00087_),
    .Q(\w[25][27] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][28]$_SDFFCE_PN0P_  (.D(_01342_),
    .DE(_00087_),
    .Q(\w[25][28] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][29]$_SDFFCE_PN0P_  (.D(_01343_),
    .DE(_00087_),
    .Q(\w[25][29] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][2]$_SDFFCE_PN0P_  (.D(_01344_),
    .DE(_00087_),
    .Q(\w[25][2] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][30]$_SDFFCE_PN0P_  (.D(_01345_),
    .DE(_00087_),
    .Q(\w[25][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][31]$_SDFFCE_PN0P_  (.D(_01346_),
    .DE(_00087_),
    .Q(\w[25][31] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][3]$_SDFFCE_PN0P_  (.D(_01347_),
    .DE(_00087_),
    .Q(\w[25][3] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][4]$_SDFFCE_PN0P_  (.D(_01348_),
    .DE(_00087_),
    .Q(\w[25][4] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][5]$_SDFFCE_PN0P_  (.D(_01349_),
    .DE(_00087_),
    .Q(\w[25][5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][6]$_SDFFCE_PN0P_  (.D(_01350_),
    .DE(_00087_),
    .Q(\w[25][6] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][7]$_SDFFCE_PN0P_  (.D(_01351_),
    .DE(_00087_),
    .Q(\w[25][7] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][8]$_SDFFCE_PN0P_  (.D(_01352_),
    .DE(_00087_),
    .Q(\w[25][8] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[25][9]$_SDFFCE_PN0P_  (.D(_01353_),
    .DE(_00087_),
    .Q(\w[25][9] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][0]$_SDFFCE_PN0P_  (.D(_01354_),
    .DE(_00118_),
    .Q(\w[26][0] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][10]$_SDFFCE_PN0P_  (.D(_01355_),
    .DE(_00118_),
    .Q(\w[26][10] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][11]$_SDFFCE_PN0P_  (.D(_01356_),
    .DE(_00118_),
    .Q(\w[26][11] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][12]$_SDFFCE_PN0P_  (.D(_01357_),
    .DE(_00118_),
    .Q(\w[26][12] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][13]$_SDFFCE_PN0P_  (.D(_01358_),
    .DE(_00118_),
    .Q(\w[26][13] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][14]$_SDFFCE_PN0P_  (.D(_01359_),
    .DE(_00118_),
    .Q(\w[26][14] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][15]$_SDFFCE_PN0P_  (.D(_01360_),
    .DE(_00118_),
    .Q(\w[26][15] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][16]$_SDFFCE_PN0P_  (.D(_01361_),
    .DE(_00118_),
    .Q(\w[26][16] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][17]$_SDFFCE_PN0P_  (.D(_01362_),
    .DE(_00118_),
    .Q(\w[26][17] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][18]$_SDFFCE_PN0P_  (.D(_01363_),
    .DE(_00118_),
    .Q(\w[26][18] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][19]$_SDFFCE_PN0P_  (.D(_01364_),
    .DE(_00118_),
    .Q(\w[26][19] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][1]$_SDFFCE_PN0P_  (.D(_01365_),
    .DE(_00118_),
    .Q(\w[26][1] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][20]$_SDFFCE_PN0P_  (.D(_01366_),
    .DE(_00118_),
    .Q(\w[26][20] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][21]$_SDFFCE_PN0P_  (.D(_01367_),
    .DE(_00118_),
    .Q(\w[26][21] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][22]$_SDFFCE_PN0P_  (.D(_01368_),
    .DE(_00118_),
    .Q(\w[26][22] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][23]$_SDFFCE_PN0P_  (.D(_01369_),
    .DE(_00118_),
    .Q(\w[26][23] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][24]$_SDFFCE_PN0P_  (.D(_01370_),
    .DE(_00118_),
    .Q(\w[26][24] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][25]$_SDFFCE_PN0P_  (.D(_01371_),
    .DE(_00118_),
    .Q(\w[26][25] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][26]$_SDFFCE_PN0P_  (.D(_01372_),
    .DE(_00118_),
    .Q(\w[26][26] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][27]$_SDFFCE_PN0P_  (.D(_01373_),
    .DE(_00118_),
    .Q(\w[26][27] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][28]$_SDFFCE_PN0P_  (.D(_01374_),
    .DE(_00118_),
    .Q(\w[26][28] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][29]$_SDFFCE_PN0P_  (.D(_01375_),
    .DE(_00118_),
    .Q(\w[26][29] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][2]$_SDFFCE_PN0P_  (.D(_01376_),
    .DE(_00118_),
    .Q(\w[26][2] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][30]$_SDFFCE_PN0P_  (.D(_01377_),
    .DE(_00118_),
    .Q(\w[26][30] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][31]$_SDFFCE_PN0P_  (.D(_01378_),
    .DE(_00118_),
    .Q(\w[26][31] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][3]$_SDFFCE_PN0P_  (.D(_01379_),
    .DE(_00118_),
    .Q(\w[26][3] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][4]$_SDFFCE_PN0P_  (.D(_01380_),
    .DE(_00118_),
    .Q(\w[26][4] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][5]$_SDFFCE_PN0P_  (.D(_01381_),
    .DE(_00118_),
    .Q(\w[26][5] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][6]$_SDFFCE_PN0P_  (.D(_01382_),
    .DE(_00118_),
    .Q(\w[26][6] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][7]$_SDFFCE_PN0P_  (.D(_01383_),
    .DE(_00118_),
    .Q(\w[26][7] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][8]$_SDFFCE_PN0P_  (.D(_01384_),
    .DE(_00118_),
    .Q(\w[26][8] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[26][9]$_SDFFCE_PN0P_  (.D(_01385_),
    .DE(_00118_),
    .Q(\w[26][9] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][0]$_SDFFCE_PN0P_  (.D(_01386_),
    .DE(_00086_),
    .Q(\w[27][0] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][10]$_SDFFCE_PN0P_  (.D(_01387_),
    .DE(_00086_),
    .Q(\w[27][10] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][11]$_SDFFCE_PN0P_  (.D(_01388_),
    .DE(_00086_),
    .Q(\w[27][11] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][12]$_SDFFCE_PN0P_  (.D(_01389_),
    .DE(_00086_),
    .Q(\w[27][12] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][13]$_SDFFCE_PN0P_  (.D(_01390_),
    .DE(_00086_),
    .Q(\w[27][13] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][14]$_SDFFCE_PN0P_  (.D(_01391_),
    .DE(_00086_),
    .Q(\w[27][14] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][15]$_SDFFCE_PN0P_  (.D(_01392_),
    .DE(_00086_),
    .Q(\w[27][15] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][16]$_SDFFCE_PN0P_  (.D(_01393_),
    .DE(_00086_),
    .Q(\w[27][16] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][17]$_SDFFCE_PN0P_  (.D(_01394_),
    .DE(_00086_),
    .Q(\w[27][17] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][18]$_SDFFCE_PN0P_  (.D(_01395_),
    .DE(_00086_),
    .Q(\w[27][18] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][19]$_SDFFCE_PN0P_  (.D(_01396_),
    .DE(_00086_),
    .Q(\w[27][19] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][1]$_SDFFCE_PN0P_  (.D(_01397_),
    .DE(_00086_),
    .Q(\w[27][1] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][20]$_SDFFCE_PN0P_  (.D(_01398_),
    .DE(_00086_),
    .Q(\w[27][20] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][21]$_SDFFCE_PN0P_  (.D(_01399_),
    .DE(_00086_),
    .Q(\w[27][21] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][22]$_SDFFCE_PN0P_  (.D(_01400_),
    .DE(_00086_),
    .Q(\w[27][22] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][23]$_SDFFCE_PN0P_  (.D(_01401_),
    .DE(_00086_),
    .Q(\w[27][23] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][24]$_SDFFCE_PN0P_  (.D(_01402_),
    .DE(_00086_),
    .Q(\w[27][24] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][25]$_SDFFCE_PN0P_  (.D(_01403_),
    .DE(_00086_),
    .Q(\w[27][25] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][26]$_SDFFCE_PN0P_  (.D(_01404_),
    .DE(_00086_),
    .Q(\w[27][26] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][27]$_SDFFCE_PN0P_  (.D(_01405_),
    .DE(_00086_),
    .Q(\w[27][27] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][28]$_SDFFCE_PN0P_  (.D(_01406_),
    .DE(_00086_),
    .Q(\w[27][28] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][29]$_SDFFCE_PN0P_  (.D(_01407_),
    .DE(_00086_),
    .Q(\w[27][29] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][2]$_SDFFCE_PN0P_  (.D(_01408_),
    .DE(_00086_),
    .Q(\w[27][2] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][30]$_SDFFCE_PN0P_  (.D(_01409_),
    .DE(_00086_),
    .Q(\w[27][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][31]$_SDFFCE_PN0P_  (.D(_01410_),
    .DE(_00086_),
    .Q(\w[27][31] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][3]$_SDFFCE_PN0P_  (.D(_01411_),
    .DE(_00086_),
    .Q(\w[27][3] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][4]$_SDFFCE_PN0P_  (.D(_01412_),
    .DE(_00086_),
    .Q(\w[27][4] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][5]$_SDFFCE_PN0P_  (.D(_01413_),
    .DE(_00086_),
    .Q(\w[27][5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][6]$_SDFFCE_PN0P_  (.D(_01414_),
    .DE(_00086_),
    .Q(\w[27][6] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][7]$_SDFFCE_PN0P_  (.D(_01415_),
    .DE(_00086_),
    .Q(\w[27][7] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][8]$_SDFFCE_PN0P_  (.D(_01416_),
    .DE(_00086_),
    .Q(\w[27][8] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[27][9]$_SDFFCE_PN0P_  (.D(_01417_),
    .DE(_00086_),
    .Q(\w[27][9] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][0]$_SDFFCE_PN0P_  (.D(_01418_),
    .DE(_00117_),
    .Q(\w[28][0] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][10]$_SDFFCE_PN0P_  (.D(_01419_),
    .DE(_00117_),
    .Q(\w[28][10] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][11]$_SDFFCE_PN0P_  (.D(_01420_),
    .DE(_00117_),
    .Q(\w[28][11] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][12]$_SDFFCE_PN0P_  (.D(_01421_),
    .DE(_00117_),
    .Q(\w[28][12] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][13]$_SDFFCE_PN0P_  (.D(_01422_),
    .DE(_00117_),
    .Q(\w[28][13] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][14]$_SDFFCE_PN0P_  (.D(_01423_),
    .DE(_00117_),
    .Q(\w[28][14] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][15]$_SDFFCE_PN0P_  (.D(_01424_),
    .DE(_00117_),
    .Q(\w[28][15] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][16]$_SDFFCE_PN0P_  (.D(_01425_),
    .DE(_00117_),
    .Q(\w[28][16] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][17]$_SDFFCE_PN0P_  (.D(_01426_),
    .DE(_00117_),
    .Q(\w[28][17] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][18]$_SDFFCE_PN0P_  (.D(_01427_),
    .DE(_00117_),
    .Q(\w[28][18] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][19]$_SDFFCE_PN0P_  (.D(_01428_),
    .DE(_00117_),
    .Q(\w[28][19] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][1]$_SDFFCE_PN0P_  (.D(_01429_),
    .DE(_00117_),
    .Q(\w[28][1] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][20]$_SDFFCE_PN0P_  (.D(_01430_),
    .DE(_00117_),
    .Q(\w[28][20] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][21]$_SDFFCE_PN0P_  (.D(_01431_),
    .DE(_00117_),
    .Q(\w[28][21] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][22]$_SDFFCE_PN0P_  (.D(_01432_),
    .DE(_00117_),
    .Q(\w[28][22] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][23]$_SDFFCE_PN0P_  (.D(_01433_),
    .DE(_00117_),
    .Q(\w[28][23] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][24]$_SDFFCE_PN0P_  (.D(_01434_),
    .DE(_00117_),
    .Q(\w[28][24] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][25]$_SDFFCE_PN0P_  (.D(_01435_),
    .DE(_00117_),
    .Q(\w[28][25] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][26]$_SDFFCE_PN0P_  (.D(_01436_),
    .DE(_00117_),
    .Q(\w[28][26] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][27]$_SDFFCE_PN0P_  (.D(_01437_),
    .DE(_00117_),
    .Q(\w[28][27] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][28]$_SDFFCE_PN0P_  (.D(_01438_),
    .DE(_00117_),
    .Q(\w[28][28] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][29]$_SDFFCE_PN0P_  (.D(_01439_),
    .DE(_00117_),
    .Q(\w[28][29] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][2]$_SDFFCE_PN0P_  (.D(_01440_),
    .DE(_00117_),
    .Q(\w[28][2] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][30]$_SDFFCE_PN0P_  (.D(_01441_),
    .DE(_00117_),
    .Q(\w[28][30] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][31]$_SDFFCE_PN0P_  (.D(_01442_),
    .DE(_00117_),
    .Q(\w[28][31] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][3]$_SDFFCE_PN0P_  (.D(_01443_),
    .DE(_00117_),
    .Q(\w[28][3] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][4]$_SDFFCE_PN0P_  (.D(_01444_),
    .DE(_00117_),
    .Q(\w[28][4] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][5]$_SDFFCE_PN0P_  (.D(_01445_),
    .DE(_00117_),
    .Q(\w[28][5] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][6]$_SDFFCE_PN0P_  (.D(_01446_),
    .DE(_00117_),
    .Q(\w[28][6] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][7]$_SDFFCE_PN0P_  (.D(_01447_),
    .DE(_00117_),
    .Q(\w[28][7] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][8]$_SDFFCE_PN0P_  (.D(_01448_),
    .DE(_00117_),
    .Q(\w[28][8] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[28][9]$_SDFFCE_PN0P_  (.D(_01449_),
    .DE(_00117_),
    .Q(\w[28][9] ),
    .CLK(clknet_leaf_137_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][0]$_SDFFCE_PN0P_  (.D(_01450_),
    .DE(_00085_),
    .Q(\w[29][0] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][10]$_SDFFCE_PN0P_  (.D(_01451_),
    .DE(_00085_),
    .Q(\w[29][10] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][11]$_SDFFCE_PN0P_  (.D(_01452_),
    .DE(_00085_),
    .Q(\w[29][11] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][12]$_SDFFCE_PN0P_  (.D(_01453_),
    .DE(_00085_),
    .Q(\w[29][12] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][13]$_SDFFCE_PN0P_  (.D(_01454_),
    .DE(_00085_),
    .Q(\w[29][13] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][14]$_SDFFCE_PN0P_  (.D(_01455_),
    .DE(_00085_),
    .Q(\w[29][14] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][15]$_SDFFCE_PN0P_  (.D(_01456_),
    .DE(_00085_),
    .Q(\w[29][15] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][16]$_SDFFCE_PN0P_  (.D(_01457_),
    .DE(_00085_),
    .Q(\w[29][16] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][17]$_SDFFCE_PN0P_  (.D(_01458_),
    .DE(_00085_),
    .Q(\w[29][17] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][18]$_SDFFCE_PN0P_  (.D(_01459_),
    .DE(_00085_),
    .Q(\w[29][18] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][19]$_SDFFCE_PN0P_  (.D(_01460_),
    .DE(_00085_),
    .Q(\w[29][19] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][1]$_SDFFCE_PN0P_  (.D(_01461_),
    .DE(_00085_),
    .Q(\w[29][1] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][20]$_SDFFCE_PN0P_  (.D(_01462_),
    .DE(_00085_),
    .Q(\w[29][20] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][21]$_SDFFCE_PN0P_  (.D(_01463_),
    .DE(_00085_),
    .Q(\w[29][21] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][22]$_SDFFCE_PN0P_  (.D(_01464_),
    .DE(_00085_),
    .Q(\w[29][22] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][23]$_SDFFCE_PN0P_  (.D(_01465_),
    .DE(_00085_),
    .Q(\w[29][23] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][24]$_SDFFCE_PN0P_  (.D(_01466_),
    .DE(_00085_),
    .Q(\w[29][24] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][25]$_SDFFCE_PN0P_  (.D(_01467_),
    .DE(_00085_),
    .Q(\w[29][25] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][26]$_SDFFCE_PN0P_  (.D(_01468_),
    .DE(_00085_),
    .Q(\w[29][26] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][27]$_SDFFCE_PN0P_  (.D(_01469_),
    .DE(_00085_),
    .Q(\w[29][27] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][28]$_SDFFCE_PN0P_  (.D(_01470_),
    .DE(_00085_),
    .Q(\w[29][28] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][29]$_SDFFCE_PN0P_  (.D(_01471_),
    .DE(_00085_),
    .Q(\w[29][29] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][2]$_SDFFCE_PN0P_  (.D(_01472_),
    .DE(_00085_),
    .Q(\w[29][2] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][30]$_SDFFCE_PN0P_  (.D(_01473_),
    .DE(_00085_),
    .Q(\w[29][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][31]$_SDFFCE_PN0P_  (.D(_01474_),
    .DE(_00085_),
    .Q(\w[29][31] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][3]$_SDFFCE_PN0P_  (.D(_01475_),
    .DE(_00085_),
    .Q(\w[29][3] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][4]$_SDFFCE_PN0P_  (.D(_01476_),
    .DE(_00085_),
    .Q(\w[29][4] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][5]$_SDFFCE_PN0P_  (.D(_01477_),
    .DE(_00085_),
    .Q(\w[29][5] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][6]$_SDFFCE_PN0P_  (.D(_01478_),
    .DE(_00085_),
    .Q(\w[29][6] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][7]$_SDFFCE_PN0P_  (.D(_01479_),
    .DE(_00085_),
    .Q(\w[29][7] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][8]$_SDFFCE_PN0P_  (.D(_01480_),
    .DE(_00085_),
    .Q(\w[29][8] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[29][9]$_SDFFCE_PN0P_  (.D(_01481_),
    .DE(_00085_),
    .Q(\w[29][9] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][0]$_DFFE_PP_  (.D(_00385_),
    .DE(_00116_),
    .Q(\w[2][0] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][10]$_DFFE_PP_  (.D(_00386_),
    .DE(_00116_),
    .Q(\w[2][10] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][11]$_DFFE_PP_  (.D(_00387_),
    .DE(_00116_),
    .Q(\w[2][11] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][12]$_DFFE_PP_  (.D(_00388_),
    .DE(_00116_),
    .Q(\w[2][12] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][13]$_DFFE_PP_  (.D(_00389_),
    .DE(_00116_),
    .Q(\w[2][13] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][14]$_DFFE_PP_  (.D(_00390_),
    .DE(_00116_),
    .Q(\w[2][14] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][15]$_DFFE_PP_  (.D(_00391_),
    .DE(_00116_),
    .Q(\w[2][15] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][16]$_DFFE_PP_  (.D(_00392_),
    .DE(_00116_),
    .Q(\w[2][16] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][17]$_DFFE_PP_  (.D(_00393_),
    .DE(_00116_),
    .Q(\w[2][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][18]$_DFFE_PP_  (.D(_00394_),
    .DE(_00116_),
    .Q(\w[2][18] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][19]$_DFFE_PP_  (.D(_00395_),
    .DE(_00116_),
    .Q(\w[2][19] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][1]$_DFFE_PP_  (.D(_00396_),
    .DE(_00116_),
    .Q(\w[2][1] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][20]$_DFFE_PP_  (.D(_00397_),
    .DE(_00116_),
    .Q(\w[2][20] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][21]$_DFFE_PP_  (.D(_00398_),
    .DE(_00116_),
    .Q(\w[2][21] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][22]$_DFFE_PP_  (.D(_00399_),
    .DE(_00116_),
    .Q(\w[2][22] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][23]$_DFFE_PP_  (.D(_00400_),
    .DE(_00116_),
    .Q(\w[2][23] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][24]$_DFFE_PP_  (.D(_00401_),
    .DE(_00116_),
    .Q(\w[2][24] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][25]$_DFFE_PP_  (.D(_00402_),
    .DE(_00116_),
    .Q(\w[2][25] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][26]$_DFFE_PP_  (.D(_00403_),
    .DE(_00116_),
    .Q(\w[2][26] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][27]$_DFFE_PP_  (.D(_00404_),
    .DE(_00116_),
    .Q(\w[2][27] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][28]$_DFFE_PP_  (.D(_00405_),
    .DE(_00116_),
    .Q(\w[2][28] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][29]$_DFFE_PP_  (.D(_00406_),
    .DE(_00116_),
    .Q(\w[2][29] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][2]$_DFFE_PP_  (.D(_00407_),
    .DE(_00116_),
    .Q(\w[2][2] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][30]$_DFFE_PP_  (.D(_00408_),
    .DE(_00116_),
    .Q(\w[2][30] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][31]$_DFFE_PP_  (.D(_00409_),
    .DE(_00116_),
    .Q(\w[2][31] ),
    .CLK(clknet_leaf_96_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][3]$_DFFE_PP_  (.D(_00410_),
    .DE(_00116_),
    .Q(\w[2][3] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][4]$_DFFE_PP_  (.D(_00411_),
    .DE(_00116_),
    .Q(\w[2][4] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][5]$_DFFE_PP_  (.D(_00412_),
    .DE(_00116_),
    .Q(\w[2][5] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][6]$_DFFE_PP_  (.D(_00413_),
    .DE(_00116_),
    .Q(\w[2][6] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][7]$_DFFE_PP_  (.D(_00414_),
    .DE(_00116_),
    .Q(\w[2][7] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][8]$_DFFE_PP_  (.D(_00415_),
    .DE(_00116_),
    .Q(\w[2][8] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[2][9]$_DFFE_PP_  (.D(_00416_),
    .DE(_00116_),
    .Q(\w[2][9] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][0]$_SDFFCE_PN0P_  (.D(_01482_),
    .DE(_00115_),
    .Q(\w[30][0] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][10]$_SDFFCE_PN0P_  (.D(_01483_),
    .DE(_00115_),
    .Q(\w[30][10] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][11]$_SDFFCE_PN0P_  (.D(_01484_),
    .DE(_00115_),
    .Q(\w[30][11] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][12]$_SDFFCE_PN0P_  (.D(_01485_),
    .DE(_00115_),
    .Q(\w[30][12] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][13]$_SDFFCE_PN0P_  (.D(_01486_),
    .DE(_00115_),
    .Q(\w[30][13] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][14]$_SDFFCE_PN0P_  (.D(_01487_),
    .DE(_00115_),
    .Q(\w[30][14] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][15]$_SDFFCE_PN0P_  (.D(_01488_),
    .DE(_00115_),
    .Q(\w[30][15] ),
    .CLK(clknet_leaf_61_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][16]$_SDFFCE_PN0P_  (.D(_01489_),
    .DE(_00115_),
    .Q(\w[30][16] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][17]$_SDFFCE_PN0P_  (.D(_01490_),
    .DE(_00115_),
    .Q(\w[30][17] ),
    .CLK(clknet_leaf_95_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][18]$_SDFFCE_PN0P_  (.D(_01491_),
    .DE(_00115_),
    .Q(\w[30][18] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][19]$_SDFFCE_PN0P_  (.D(_01492_),
    .DE(_00115_),
    .Q(\w[30][19] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][1]$_SDFFCE_PN0P_  (.D(_01493_),
    .DE(_00115_),
    .Q(\w[30][1] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][20]$_SDFFCE_PN0P_  (.D(_01494_),
    .DE(_00115_),
    .Q(\w[30][20] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][21]$_SDFFCE_PN0P_  (.D(_01495_),
    .DE(_00115_),
    .Q(\w[30][21] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][22]$_SDFFCE_PN0P_  (.D(_01496_),
    .DE(_00115_),
    .Q(\w[30][22] ),
    .CLK(clknet_leaf_144_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][23]$_SDFFCE_PN0P_  (.D(_01497_),
    .DE(_00115_),
    .Q(\w[30][23] ),
    .CLK(clknet_leaf_90_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][24]$_SDFFCE_PN0P_  (.D(_01498_),
    .DE(_00115_),
    .Q(\w[30][24] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][25]$_SDFFCE_PN0P_  (.D(_01499_),
    .DE(_00115_),
    .Q(\w[30][25] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][26]$_SDFFCE_PN0P_  (.D(_01500_),
    .DE(_00115_),
    .Q(\w[30][26] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][27]$_SDFFCE_PN0P_  (.D(_01501_),
    .DE(_00115_),
    .Q(\w[30][27] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][28]$_SDFFCE_PN0P_  (.D(_01502_),
    .DE(_00115_),
    .Q(\w[30][28] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][29]$_SDFFCE_PN0P_  (.D(_01503_),
    .DE(_00115_),
    .Q(\w[30][29] ),
    .CLK(clknet_leaf_78_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][2]$_SDFFCE_PN0P_  (.D(_01504_),
    .DE(_00115_),
    .Q(\w[30][2] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][30]$_SDFFCE_PN0P_  (.D(_01505_),
    .DE(_00115_),
    .Q(\w[30][30] ),
    .CLK(clknet_leaf_75_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][31]$_SDFFCE_PN0P_  (.D(_01506_),
    .DE(_00115_),
    .Q(\w[30][31] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][3]$_SDFFCE_PN0P_  (.D(_01507_),
    .DE(_00115_),
    .Q(\w[30][3] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][4]$_SDFFCE_PN0P_  (.D(_01508_),
    .DE(_00115_),
    .Q(\w[30][4] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][5]$_SDFFCE_PN0P_  (.D(_01509_),
    .DE(_00115_),
    .Q(\w[30][5] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][6]$_SDFFCE_PN0P_  (.D(_01510_),
    .DE(_00115_),
    .Q(\w[30][6] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][7]$_SDFFCE_PN0P_  (.D(_01511_),
    .DE(_00115_),
    .Q(\w[30][7] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][8]$_SDFFCE_PN0P_  (.D(_01512_),
    .DE(_00115_),
    .Q(\w[30][8] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[30][9]$_SDFFCE_PN0P_  (.D(_01513_),
    .DE(_00115_),
    .Q(\w[30][9] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][0]$_SDFFCE_PN0P_  (.D(_01514_),
    .DE(_00084_),
    .Q(\w[31][0] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][10]$_SDFFCE_PN0P_  (.D(_01515_),
    .DE(_00084_),
    .Q(\w[31][10] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][11]$_SDFFCE_PN0P_  (.D(_01516_),
    .DE(_00084_),
    .Q(\w[31][11] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][12]$_SDFFCE_PN0P_  (.D(_01517_),
    .DE(_00084_),
    .Q(\w[31][12] ),
    .CLK(clknet_leaf_225_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][13]$_SDFFCE_PN0P_  (.D(_01518_),
    .DE(_00084_),
    .Q(\w[31][13] ),
    .CLK(clknet_leaf_242_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][14]$_SDFFCE_PN0P_  (.D(_01519_),
    .DE(_00084_),
    .Q(\w[31][14] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][15]$_SDFFCE_PN0P_  (.D(_01520_),
    .DE(_00084_),
    .Q(\w[31][15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][16]$_SDFFCE_PN0P_  (.D(_01521_),
    .DE(_00084_),
    .Q(\w[31][16] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][17]$_SDFFCE_PN0P_  (.D(_01522_),
    .DE(_00084_),
    .Q(\w[31][17] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][18]$_SDFFCE_PN0P_  (.D(_01523_),
    .DE(_00084_),
    .Q(\w[31][18] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][19]$_SDFFCE_PN0P_  (.D(_01524_),
    .DE(_00084_),
    .Q(\w[31][19] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][1]$_SDFFCE_PN0P_  (.D(_01525_),
    .DE(_00084_),
    .Q(\w[31][1] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][20]$_SDFFCE_PN0P_  (.D(_01526_),
    .DE(_00084_),
    .Q(\w[31][20] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][21]$_SDFFCE_PN0P_  (.D(_01527_),
    .DE(_00084_),
    .Q(\w[31][21] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][22]$_SDFFCE_PN0P_  (.D(_01528_),
    .DE(_00084_),
    .Q(\w[31][22] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][23]$_SDFFCE_PN0P_  (.D(_01529_),
    .DE(_00084_),
    .Q(\w[31][23] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][24]$_SDFFCE_PN0P_  (.D(_01530_),
    .DE(_00084_),
    .Q(\w[31][24] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][25]$_SDFFCE_PN0P_  (.D(_01531_),
    .DE(_00084_),
    .Q(\w[31][25] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][26]$_SDFFCE_PN0P_  (.D(_01532_),
    .DE(_00084_),
    .Q(\w[31][26] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][27]$_SDFFCE_PN0P_  (.D(_01533_),
    .DE(_00084_),
    .Q(\w[31][27] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][28]$_SDFFCE_PN0P_  (.D(_01534_),
    .DE(_00084_),
    .Q(\w[31][28] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][29]$_SDFFCE_PN0P_  (.D(_01535_),
    .DE(_00084_),
    .Q(\w[31][29] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][2]$_SDFFCE_PN0P_  (.D(_01536_),
    .DE(_00084_),
    .Q(\w[31][2] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][30]$_SDFFCE_PN0P_  (.D(_01537_),
    .DE(_00084_),
    .Q(\w[31][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][31]$_SDFFCE_PN0P_  (.D(_01538_),
    .DE(_00084_),
    .Q(\w[31][31] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][3]$_SDFFCE_PN0P_  (.D(_01539_),
    .DE(_00084_),
    .Q(\w[31][3] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][4]$_SDFFCE_PN0P_  (.D(_01540_),
    .DE(_00084_),
    .Q(\w[31][4] ),
    .CLK(clknet_leaf_274_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][5]$_SDFFCE_PN0P_  (.D(_01541_),
    .DE(_00084_),
    .Q(\w[31][5] ),
    .CLK(clknet_leaf_1_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][6]$_SDFFCE_PN0P_  (.D(_01542_),
    .DE(_00084_),
    .Q(\w[31][6] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][7]$_SDFFCE_PN0P_  (.D(_01543_),
    .DE(_00084_),
    .Q(\w[31][7] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][8]$_SDFFCE_PN0P_  (.D(_01544_),
    .DE(_00084_),
    .Q(\w[31][8] ),
    .CLK(clknet_leaf_265_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[31][9]$_SDFFCE_PN0P_  (.D(_01545_),
    .DE(_00084_),
    .Q(\w[31][9] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][0]$_SDFFCE_PN0P_  (.D(_01546_),
    .DE(_00114_),
    .Q(\w[32][0] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][10]$_SDFFCE_PN0P_  (.D(_01547_),
    .DE(_00114_),
    .Q(\w[32][10] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][11]$_SDFFCE_PN0P_  (.D(_01548_),
    .DE(_00114_),
    .Q(\w[32][11] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][12]$_SDFFCE_PN0P_  (.D(_01549_),
    .DE(_00114_),
    .Q(\w[32][12] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][13]$_SDFFCE_PN0P_  (.D(_01550_),
    .DE(_00114_),
    .Q(\w[32][13] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][14]$_SDFFCE_PN0P_  (.D(_01551_),
    .DE(_00114_),
    .Q(\w[32][14] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][15]$_SDFFCE_PN0P_  (.D(_01552_),
    .DE(_00114_),
    .Q(\w[32][15] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][16]$_SDFFCE_PN0P_  (.D(_01553_),
    .DE(_00114_),
    .Q(\w[32][16] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][17]$_SDFFCE_PN0P_  (.D(_01554_),
    .DE(_00114_),
    .Q(\w[32][17] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][18]$_SDFFCE_PN0P_  (.D(_01555_),
    .DE(_00114_),
    .Q(\w[32][18] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][19]$_SDFFCE_PN0P_  (.D(_01556_),
    .DE(_00114_),
    .Q(\w[32][19] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][1]$_SDFFCE_PN0P_  (.D(_01557_),
    .DE(_00114_),
    .Q(\w[32][1] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][20]$_SDFFCE_PN0P_  (.D(_01558_),
    .DE(_00114_),
    .Q(\w[32][20] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][21]$_SDFFCE_PN0P_  (.D(_01559_),
    .DE(_00114_),
    .Q(\w[32][21] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][22]$_SDFFCE_PN0P_  (.D(_01560_),
    .DE(_00114_),
    .Q(\w[32][22] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][23]$_SDFFCE_PN0P_  (.D(_01561_),
    .DE(_00114_),
    .Q(\w[32][23] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][24]$_SDFFCE_PN0P_  (.D(_01562_),
    .DE(_00114_),
    .Q(\w[32][24] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][25]$_SDFFCE_PN0P_  (.D(_01563_),
    .DE(_00114_),
    .Q(\w[32][25] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][26]$_SDFFCE_PN0P_  (.D(_01564_),
    .DE(_00114_),
    .Q(\w[32][26] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][27]$_SDFFCE_PN0P_  (.D(_01565_),
    .DE(_00114_),
    .Q(\w[32][27] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][28]$_SDFFCE_PN0P_  (.D(_01566_),
    .DE(_00114_),
    .Q(\w[32][28] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][29]$_SDFFCE_PN0P_  (.D(_01567_),
    .DE(_00114_),
    .Q(\w[32][29] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][2]$_SDFFCE_PN0P_  (.D(_01568_),
    .DE(_00114_),
    .Q(\w[32][2] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][30]$_SDFFCE_PN0P_  (.D(_01569_),
    .DE(_00114_),
    .Q(\w[32][30] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][31]$_SDFFCE_PN0P_  (.D(_01570_),
    .DE(_00114_),
    .Q(\w[32][31] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][3]$_SDFFCE_PN0P_  (.D(_01571_),
    .DE(_00114_),
    .Q(\w[32][3] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][4]$_SDFFCE_PN0P_  (.D(_01572_),
    .DE(_00114_),
    .Q(\w[32][4] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][5]$_SDFFCE_PN0P_  (.D(_01573_),
    .DE(_00114_),
    .Q(\w[32][5] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][6]$_SDFFCE_PN0P_  (.D(_01574_),
    .DE(_00114_),
    .Q(\w[32][6] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][7]$_SDFFCE_PN0P_  (.D(_01575_),
    .DE(_00114_),
    .Q(\w[32][7] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][8]$_SDFFCE_PN0P_  (.D(_01576_),
    .DE(_00114_),
    .Q(\w[32][8] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[32][9]$_SDFFCE_PN0P_  (.D(_01577_),
    .DE(_00114_),
    .Q(\w[32][9] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][0]$_SDFFCE_PN0P_  (.D(_01578_),
    .DE(_00083_),
    .Q(\w[33][0] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][10]$_SDFFCE_PN0P_  (.D(_01579_),
    .DE(_00083_),
    .Q(\w[33][10] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][11]$_SDFFCE_PN0P_  (.D(_01580_),
    .DE(_00083_),
    .Q(\w[33][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][12]$_SDFFCE_PN0P_  (.D(_01581_),
    .DE(_00083_),
    .Q(\w[33][12] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][13]$_SDFFCE_PN0P_  (.D(_01582_),
    .DE(_00083_),
    .Q(\w[33][13] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][14]$_SDFFCE_PN0P_  (.D(_01583_),
    .DE(_00083_),
    .Q(\w[33][14] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][15]$_SDFFCE_PN0P_  (.D(_01584_),
    .DE(_00083_),
    .Q(\w[33][15] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][16]$_SDFFCE_PN0P_  (.D(_01585_),
    .DE(_00083_),
    .Q(\w[33][16] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][17]$_SDFFCE_PN0P_  (.D(_01586_),
    .DE(_00083_),
    .Q(\w[33][17] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][18]$_SDFFCE_PN0P_  (.D(_01587_),
    .DE(_00083_),
    .Q(\w[33][18] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][19]$_SDFFCE_PN0P_  (.D(_01588_),
    .DE(_00083_),
    .Q(\w[33][19] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][1]$_SDFFCE_PN0P_  (.D(_01589_),
    .DE(_00083_),
    .Q(\w[33][1] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][20]$_SDFFCE_PN0P_  (.D(_01590_),
    .DE(_00083_),
    .Q(\w[33][20] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][21]$_SDFFCE_PN0P_  (.D(_01591_),
    .DE(_00083_),
    .Q(\w[33][21] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][22]$_SDFFCE_PN0P_  (.D(_01592_),
    .DE(_00083_),
    .Q(\w[33][22] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][23]$_SDFFCE_PN0P_  (.D(_01593_),
    .DE(_00083_),
    .Q(\w[33][23] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][24]$_SDFFCE_PN0P_  (.D(_01594_),
    .DE(_00083_),
    .Q(\w[33][24] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][25]$_SDFFCE_PN0P_  (.D(_01595_),
    .DE(_00083_),
    .Q(\w[33][25] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][26]$_SDFFCE_PN0P_  (.D(_01596_),
    .DE(_00083_),
    .Q(\w[33][26] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][27]$_SDFFCE_PN0P_  (.D(_01597_),
    .DE(_00083_),
    .Q(\w[33][27] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][28]$_SDFFCE_PN0P_  (.D(_01598_),
    .DE(_00083_),
    .Q(\w[33][28] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][29]$_SDFFCE_PN0P_  (.D(_01599_),
    .DE(_00083_),
    .Q(\w[33][29] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][2]$_SDFFCE_PN0P_  (.D(_01600_),
    .DE(_00083_),
    .Q(\w[33][2] ),
    .CLK(clknet_leaf_275_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][30]$_SDFFCE_PN0P_  (.D(_01601_),
    .DE(_00083_),
    .Q(\w[33][30] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][31]$_SDFFCE_PN0P_  (.D(_01602_),
    .DE(_00083_),
    .Q(\w[33][31] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][3]$_SDFFCE_PN0P_  (.D(_01603_),
    .DE(_00083_),
    .Q(\w[33][3] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][4]$_SDFFCE_PN0P_  (.D(_01604_),
    .DE(_00083_),
    .Q(\w[33][4] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][5]$_SDFFCE_PN0P_  (.D(_01605_),
    .DE(_00083_),
    .Q(\w[33][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][6]$_SDFFCE_PN0P_  (.D(_01606_),
    .DE(_00083_),
    .Q(\w[33][6] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][7]$_SDFFCE_PN0P_  (.D(_01607_),
    .DE(_00083_),
    .Q(\w[33][7] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][8]$_SDFFCE_PN0P_  (.D(_01608_),
    .DE(_00083_),
    .Q(\w[33][8] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[33][9]$_SDFFCE_PN0P_  (.D(_01609_),
    .DE(_00083_),
    .Q(\w[33][9] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][0]$_SDFFCE_PN0P_  (.D(_01610_),
    .DE(_00113_),
    .Q(\w[34][0] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][10]$_SDFFCE_PN0P_  (.D(_01611_),
    .DE(_00113_),
    .Q(\w[34][10] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][11]$_SDFFCE_PN0P_  (.D(_01612_),
    .DE(_00113_),
    .Q(\w[34][11] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][12]$_SDFFCE_PN0P_  (.D(_01613_),
    .DE(_00113_),
    .Q(\w[34][12] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][13]$_SDFFCE_PN0P_  (.D(_01614_),
    .DE(_00113_),
    .Q(\w[34][13] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][14]$_SDFFCE_PN0P_  (.D(_01615_),
    .DE(_00113_),
    .Q(\w[34][14] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][15]$_SDFFCE_PN0P_  (.D(_01616_),
    .DE(_00113_),
    .Q(\w[34][15] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][16]$_SDFFCE_PN0P_  (.D(_01617_),
    .DE(_00113_),
    .Q(\w[34][16] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][17]$_SDFFCE_PN0P_  (.D(_01618_),
    .DE(_00113_),
    .Q(\w[34][17] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][18]$_SDFFCE_PN0P_  (.D(_01619_),
    .DE(_00113_),
    .Q(\w[34][18] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][19]$_SDFFCE_PN0P_  (.D(_01620_),
    .DE(_00113_),
    .Q(\w[34][19] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][1]$_SDFFCE_PN0P_  (.D(_01621_),
    .DE(_00113_),
    .Q(\w[34][1] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][20]$_SDFFCE_PN0P_  (.D(_01622_),
    .DE(_00113_),
    .Q(\w[34][20] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][21]$_SDFFCE_PN0P_  (.D(_01623_),
    .DE(_00113_),
    .Q(\w[34][21] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][22]$_SDFFCE_PN0P_  (.D(_01624_),
    .DE(_00113_),
    .Q(\w[34][22] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][23]$_SDFFCE_PN0P_  (.D(_01625_),
    .DE(_00113_),
    .Q(\w[34][23] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][24]$_SDFFCE_PN0P_  (.D(_01626_),
    .DE(_00113_),
    .Q(\w[34][24] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][25]$_SDFFCE_PN0P_  (.D(_01627_),
    .DE(_00113_),
    .Q(\w[34][25] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][26]$_SDFFCE_PN0P_  (.D(_01628_),
    .DE(_00113_),
    .Q(\w[34][26] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][27]$_SDFFCE_PN0P_  (.D(_01629_),
    .DE(_00113_),
    .Q(\w[34][27] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][28]$_SDFFCE_PN0P_  (.D(_01630_),
    .DE(_00113_),
    .Q(\w[34][28] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][29]$_SDFFCE_PN0P_  (.D(_01631_),
    .DE(_00113_),
    .Q(\w[34][29] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][2]$_SDFFCE_PN0P_  (.D(_01632_),
    .DE(_00113_),
    .Q(\w[34][2] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][30]$_SDFFCE_PN0P_  (.D(_01633_),
    .DE(_00113_),
    .Q(\w[34][30] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][31]$_SDFFCE_PN0P_  (.D(_01634_),
    .DE(_00113_),
    .Q(\w[34][31] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][3]$_SDFFCE_PN0P_  (.D(_01635_),
    .DE(_00113_),
    .Q(\w[34][3] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][4]$_SDFFCE_PN0P_  (.D(_01636_),
    .DE(_00113_),
    .Q(\w[34][4] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][5]$_SDFFCE_PN0P_  (.D(_01637_),
    .DE(_00113_),
    .Q(\w[34][5] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][6]$_SDFFCE_PN0P_  (.D(_01638_),
    .DE(_00113_),
    .Q(\w[34][6] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][7]$_SDFFCE_PN0P_  (.D(_01639_),
    .DE(_00113_),
    .Q(\w[34][7] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][8]$_SDFFCE_PN0P_  (.D(_01640_),
    .DE(_00113_),
    .Q(\w[34][8] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[34][9]$_SDFFCE_PN0P_  (.D(_01641_),
    .DE(_00113_),
    .Q(\w[34][9] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][0]$_SDFFCE_PN0P_  (.D(_01642_),
    .DE(_00082_),
    .Q(\w[35][0] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][10]$_SDFFCE_PN0P_  (.D(_01643_),
    .DE(_00082_),
    .Q(\w[35][10] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][11]$_SDFFCE_PN0P_  (.D(_01644_),
    .DE(_00082_),
    .Q(\w[35][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][12]$_SDFFCE_PN0P_  (.D(_01645_),
    .DE(_00082_),
    .Q(\w[35][12] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][13]$_SDFFCE_PN0P_  (.D(_01646_),
    .DE(_00082_),
    .Q(\w[35][13] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][14]$_SDFFCE_PN0P_  (.D(_01647_),
    .DE(_00082_),
    .Q(\w[35][14] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][15]$_SDFFCE_PN0P_  (.D(_01648_),
    .DE(_00082_),
    .Q(\w[35][15] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][16]$_SDFFCE_PN0P_  (.D(_01649_),
    .DE(_00082_),
    .Q(\w[35][16] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][17]$_SDFFCE_PN0P_  (.D(_01650_),
    .DE(_00082_),
    .Q(\w[35][17] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][18]$_SDFFCE_PN0P_  (.D(_01651_),
    .DE(_00082_),
    .Q(\w[35][18] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][19]$_SDFFCE_PN0P_  (.D(_01652_),
    .DE(_00082_),
    .Q(\w[35][19] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][1]$_SDFFCE_PN0P_  (.D(_01653_),
    .DE(_00082_),
    .Q(\w[35][1] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][20]$_SDFFCE_PN0P_  (.D(_01654_),
    .DE(_00082_),
    .Q(\w[35][20] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][21]$_SDFFCE_PN0P_  (.D(_01655_),
    .DE(_00082_),
    .Q(\w[35][21] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][22]$_SDFFCE_PN0P_  (.D(_01656_),
    .DE(_00082_),
    .Q(\w[35][22] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][23]$_SDFFCE_PN0P_  (.D(_01657_),
    .DE(_00082_),
    .Q(\w[35][23] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][24]$_SDFFCE_PN0P_  (.D(_01658_),
    .DE(_00082_),
    .Q(\w[35][24] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][25]$_SDFFCE_PN0P_  (.D(_01659_),
    .DE(_00082_),
    .Q(\w[35][25] ),
    .CLK(clknet_leaf_264_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][26]$_SDFFCE_PN0P_  (.D(_01660_),
    .DE(_00082_),
    .Q(\w[35][26] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][27]$_SDFFCE_PN0P_  (.D(_01661_),
    .DE(_00082_),
    .Q(\w[35][27] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][28]$_SDFFCE_PN0P_  (.D(_01662_),
    .DE(_00082_),
    .Q(\w[35][28] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][29]$_SDFFCE_PN0P_  (.D(_01663_),
    .DE(_00082_),
    .Q(\w[35][29] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][2]$_SDFFCE_PN0P_  (.D(_01664_),
    .DE(_00082_),
    .Q(\w[35][2] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][30]$_SDFFCE_PN0P_  (.D(_01665_),
    .DE(_00082_),
    .Q(\w[35][30] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][31]$_SDFFCE_PN0P_  (.D(_01666_),
    .DE(_00082_),
    .Q(\w[35][31] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][3]$_SDFFCE_PN0P_  (.D(_01667_),
    .DE(_00082_),
    .Q(\w[35][3] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][4]$_SDFFCE_PN0P_  (.D(_01668_),
    .DE(_00082_),
    .Q(\w[35][4] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][5]$_SDFFCE_PN0P_  (.D(_01669_),
    .DE(_00082_),
    .Q(\w[35][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][6]$_SDFFCE_PN0P_  (.D(_01670_),
    .DE(_00082_),
    .Q(\w[35][6] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][7]$_SDFFCE_PN0P_  (.D(_01671_),
    .DE(_00082_),
    .Q(\w[35][7] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][8]$_SDFFCE_PN0P_  (.D(_01672_),
    .DE(_00082_),
    .Q(\w[35][8] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[35][9]$_SDFFCE_PN0P_  (.D(_01673_),
    .DE(_00082_),
    .Q(\w[35][9] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][0]$_SDFFCE_PN0P_  (.D(_01674_),
    .DE(_00112_),
    .Q(\w[36][0] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][10]$_SDFFCE_PN0P_  (.D(_01675_),
    .DE(_00112_),
    .Q(\w[36][10] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][11]$_SDFFCE_PN0P_  (.D(_01676_),
    .DE(_00112_),
    .Q(\w[36][11] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][12]$_SDFFCE_PN0P_  (.D(_01677_),
    .DE(_00112_),
    .Q(\w[36][12] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][13]$_SDFFCE_PN0P_  (.D(_01678_),
    .DE(_00112_),
    .Q(\w[36][13] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][14]$_SDFFCE_PN0P_  (.D(_01679_),
    .DE(_00112_),
    .Q(\w[36][14] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][15]$_SDFFCE_PN0P_  (.D(_01680_),
    .DE(_00112_),
    .Q(\w[36][15] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][16]$_SDFFCE_PN0P_  (.D(_01681_),
    .DE(_00112_),
    .Q(\w[36][16] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][17]$_SDFFCE_PN0P_  (.D(_01682_),
    .DE(_00112_),
    .Q(\w[36][17] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][18]$_SDFFCE_PN0P_  (.D(_01683_),
    .DE(_00112_),
    .Q(\w[36][18] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][19]$_SDFFCE_PN0P_  (.D(_01684_),
    .DE(_00112_),
    .Q(\w[36][19] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][1]$_SDFFCE_PN0P_  (.D(_01685_),
    .DE(_00112_),
    .Q(\w[36][1] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][20]$_SDFFCE_PN0P_  (.D(_01686_),
    .DE(_00112_),
    .Q(\w[36][20] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][21]$_SDFFCE_PN0P_  (.D(_01687_),
    .DE(_00112_),
    .Q(\w[36][21] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][22]$_SDFFCE_PN0P_  (.D(_01688_),
    .DE(_00112_),
    .Q(\w[36][22] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][23]$_SDFFCE_PN0P_  (.D(_01689_),
    .DE(_00112_),
    .Q(\w[36][23] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][24]$_SDFFCE_PN0P_  (.D(_01690_),
    .DE(_00112_),
    .Q(\w[36][24] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][25]$_SDFFCE_PN0P_  (.D(_01691_),
    .DE(_00112_),
    .Q(\w[36][25] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][26]$_SDFFCE_PN0P_  (.D(_01692_),
    .DE(_00112_),
    .Q(\w[36][26] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][27]$_SDFFCE_PN0P_  (.D(_01693_),
    .DE(_00112_),
    .Q(\w[36][27] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][28]$_SDFFCE_PN0P_  (.D(_01694_),
    .DE(_00112_),
    .Q(\w[36][28] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][29]$_SDFFCE_PN0P_  (.D(_01695_),
    .DE(_00112_),
    .Q(\w[36][29] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][2]$_SDFFCE_PN0P_  (.D(_01696_),
    .DE(_00112_),
    .Q(\w[36][2] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][30]$_SDFFCE_PN0P_  (.D(_01697_),
    .DE(_00112_),
    .Q(\w[36][30] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][31]$_SDFFCE_PN0P_  (.D(_01698_),
    .DE(_00112_),
    .Q(\w[36][31] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][3]$_SDFFCE_PN0P_  (.D(_01699_),
    .DE(_00112_),
    .Q(\w[36][3] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][4]$_SDFFCE_PN0P_  (.D(_01700_),
    .DE(_00112_),
    .Q(\w[36][4] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][5]$_SDFFCE_PN0P_  (.D(_01701_),
    .DE(_00112_),
    .Q(\w[36][5] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][6]$_SDFFCE_PN0P_  (.D(_01702_),
    .DE(_00112_),
    .Q(\w[36][6] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][7]$_SDFFCE_PN0P_  (.D(_01703_),
    .DE(_00112_),
    .Q(\w[36][7] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][8]$_SDFFCE_PN0P_  (.D(_01704_),
    .DE(_00112_),
    .Q(\w[36][8] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[36][9]$_SDFFCE_PN0P_  (.D(_01705_),
    .DE(_00112_),
    .Q(\w[36][9] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][0]$_SDFFCE_PN0P_  (.D(_01706_),
    .DE(_00081_),
    .Q(\w[37][0] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][10]$_SDFFCE_PN0P_  (.D(_01707_),
    .DE(_00081_),
    .Q(\w[37][10] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][11]$_SDFFCE_PN0P_  (.D(_01708_),
    .DE(_00081_),
    .Q(\w[37][11] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][12]$_SDFFCE_PN0P_  (.D(_01709_),
    .DE(_00081_),
    .Q(\w[37][12] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][13]$_SDFFCE_PN0P_  (.D(_01710_),
    .DE(_00081_),
    .Q(\w[37][13] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][14]$_SDFFCE_PN0P_  (.D(_01711_),
    .DE(_00081_),
    .Q(\w[37][14] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][15]$_SDFFCE_PN0P_  (.D(_01712_),
    .DE(_00081_),
    .Q(\w[37][15] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][16]$_SDFFCE_PN0P_  (.D(_01713_),
    .DE(_00081_),
    .Q(\w[37][16] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][17]$_SDFFCE_PN0P_  (.D(_01714_),
    .DE(_00081_),
    .Q(\w[37][17] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][18]$_SDFFCE_PN0P_  (.D(_01715_),
    .DE(_00081_),
    .Q(\w[37][18] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][19]$_SDFFCE_PN0P_  (.D(_01716_),
    .DE(_00081_),
    .Q(\w[37][19] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][1]$_SDFFCE_PN0P_  (.D(_01717_),
    .DE(_00081_),
    .Q(\w[37][1] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][20]$_SDFFCE_PN0P_  (.D(_01718_),
    .DE(_00081_),
    .Q(\w[37][20] ),
    .CLK(clknet_leaf_180_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][21]$_SDFFCE_PN0P_  (.D(_01719_),
    .DE(_00081_),
    .Q(\w[37][21] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][22]$_SDFFCE_PN0P_  (.D(_01720_),
    .DE(_00081_),
    .Q(\w[37][22] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][23]$_SDFFCE_PN0P_  (.D(_01721_),
    .DE(_00081_),
    .Q(\w[37][23] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][24]$_SDFFCE_PN0P_  (.D(_01722_),
    .DE(_00081_),
    .Q(\w[37][24] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][25]$_SDFFCE_PN0P_  (.D(_01723_),
    .DE(_00081_),
    .Q(\w[37][25] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][26]$_SDFFCE_PN0P_  (.D(_01724_),
    .DE(_00081_),
    .Q(\w[37][26] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][27]$_SDFFCE_PN0P_  (.D(_01725_),
    .DE(_00081_),
    .Q(\w[37][27] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][28]$_SDFFCE_PN0P_  (.D(_01726_),
    .DE(_00081_),
    .Q(\w[37][28] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][29]$_SDFFCE_PN0P_  (.D(_01727_),
    .DE(_00081_),
    .Q(\w[37][29] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][2]$_SDFFCE_PN0P_  (.D(_01728_),
    .DE(_00081_),
    .Q(\w[37][2] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][30]$_SDFFCE_PN0P_  (.D(_01729_),
    .DE(_00081_),
    .Q(\w[37][30] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][31]$_SDFFCE_PN0P_  (.D(_01730_),
    .DE(_00081_),
    .Q(\w[37][31] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][3]$_SDFFCE_PN0P_  (.D(_01731_),
    .DE(_00081_),
    .Q(\w[37][3] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][4]$_SDFFCE_PN0P_  (.D(_01732_),
    .DE(_00081_),
    .Q(\w[37][4] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][5]$_SDFFCE_PN0P_  (.D(_01733_),
    .DE(_00081_),
    .Q(\w[37][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][6]$_SDFFCE_PN0P_  (.D(_01734_),
    .DE(_00081_),
    .Q(\w[37][6] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][7]$_SDFFCE_PN0P_  (.D(_01735_),
    .DE(_00081_),
    .Q(\w[37][7] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][8]$_SDFFCE_PN0P_  (.D(_01736_),
    .DE(_00081_),
    .Q(\w[37][8] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[37][9]$_SDFFCE_PN0P_  (.D(_01737_),
    .DE(_00081_),
    .Q(\w[37][9] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][0]$_SDFFCE_PN0P_  (.D(_01738_),
    .DE(_00111_),
    .Q(\w[38][0] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][10]$_SDFFCE_PN0P_  (.D(_01739_),
    .DE(_00111_),
    .Q(\w[38][10] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][11]$_SDFFCE_PN0P_  (.D(_01740_),
    .DE(_00111_),
    .Q(\w[38][11] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][12]$_SDFFCE_PN0P_  (.D(_01741_),
    .DE(_00111_),
    .Q(\w[38][12] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][13]$_SDFFCE_PN0P_  (.D(_01742_),
    .DE(_00111_),
    .Q(\w[38][13] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][14]$_SDFFCE_PN0P_  (.D(_01743_),
    .DE(_00111_),
    .Q(\w[38][14] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][15]$_SDFFCE_PN0P_  (.D(_01744_),
    .DE(_00111_),
    .Q(\w[38][15] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][16]$_SDFFCE_PN0P_  (.D(_01745_),
    .DE(_00111_),
    .Q(\w[38][16] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][17]$_SDFFCE_PN0P_  (.D(_01746_),
    .DE(_00111_),
    .Q(\w[38][17] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][18]$_SDFFCE_PN0P_  (.D(_01747_),
    .DE(_00111_),
    .Q(\w[38][18] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][19]$_SDFFCE_PN0P_  (.D(_01748_),
    .DE(_00111_),
    .Q(\w[38][19] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][1]$_SDFFCE_PN0P_  (.D(_01749_),
    .DE(_00111_),
    .Q(\w[38][1] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][20]$_SDFFCE_PN0P_  (.D(_01750_),
    .DE(_00111_),
    .Q(\w[38][20] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][21]$_SDFFCE_PN0P_  (.D(_01751_),
    .DE(_00111_),
    .Q(\w[38][21] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][22]$_SDFFCE_PN0P_  (.D(_01752_),
    .DE(_00111_),
    .Q(\w[38][22] ),
    .CLK(clknet_leaf_138_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][23]$_SDFFCE_PN0P_  (.D(_01753_),
    .DE(_00111_),
    .Q(\w[38][23] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][24]$_SDFFCE_PN0P_  (.D(_01754_),
    .DE(_00111_),
    .Q(\w[38][24] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][25]$_SDFFCE_PN0P_  (.D(_01755_),
    .DE(_00111_),
    .Q(\w[38][25] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][26]$_SDFFCE_PN0P_  (.D(_01756_),
    .DE(_00111_),
    .Q(\w[38][26] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][27]$_SDFFCE_PN0P_  (.D(_01757_),
    .DE(_00111_),
    .Q(\w[38][27] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][28]$_SDFFCE_PN0P_  (.D(_01758_),
    .DE(_00111_),
    .Q(\w[38][28] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][29]$_SDFFCE_PN0P_  (.D(_01759_),
    .DE(_00111_),
    .Q(\w[38][29] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][2]$_SDFFCE_PN0P_  (.D(_01760_),
    .DE(_00111_),
    .Q(\w[38][2] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][30]$_SDFFCE_PN0P_  (.D(_01761_),
    .DE(_00111_),
    .Q(\w[38][30] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][31]$_SDFFCE_PN0P_  (.D(_01762_),
    .DE(_00111_),
    .Q(\w[38][31] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][3]$_SDFFCE_PN0P_  (.D(_01763_),
    .DE(_00111_),
    .Q(\w[38][3] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][4]$_SDFFCE_PN0P_  (.D(_01764_),
    .DE(_00111_),
    .Q(\w[38][4] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][5]$_SDFFCE_PN0P_  (.D(_01765_),
    .DE(_00111_),
    .Q(\w[38][5] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][6]$_SDFFCE_PN0P_  (.D(_01766_),
    .DE(_00111_),
    .Q(\w[38][6] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][7]$_SDFFCE_PN0P_  (.D(_01767_),
    .DE(_00111_),
    .Q(\w[38][7] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][8]$_SDFFCE_PN0P_  (.D(_01768_),
    .DE(_00111_),
    .Q(\w[38][8] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[38][9]$_SDFFCE_PN0P_  (.D(_01769_),
    .DE(_00111_),
    .Q(\w[38][9] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][0]$_SDFFCE_PN0P_  (.D(_01770_),
    .DE(net298),
    .Q(\w[39][0] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][10]$_SDFFCE_PN0P_  (.D(_01771_),
    .DE(net299),
    .Q(\w[39][10] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][11]$_SDFFCE_PN0P_  (.D(_01772_),
    .DE(_00080_),
    .Q(\w[39][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][12]$_SDFFCE_PN0P_  (.D(_01773_),
    .DE(net299),
    .Q(\w[39][12] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][13]$_SDFFCE_PN0P_  (.D(_01774_),
    .DE(_00080_),
    .Q(\w[39][13] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][14]$_SDFFCE_PN0P_  (.D(_01775_),
    .DE(net298),
    .Q(\w[39][14] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][15]$_SDFFCE_PN0P_  (.D(_01776_),
    .DE(_00080_),
    .Q(\w[39][15] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][16]$_SDFFCE_PN0P_  (.D(_01777_),
    .DE(net299),
    .Q(\w[39][16] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][17]$_SDFFCE_PN0P_  (.D(_01778_),
    .DE(net298),
    .Q(\w[39][17] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][18]$_SDFFCE_PN0P_  (.D(_01779_),
    .DE(net299),
    .Q(\w[39][18] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][19]$_SDFFCE_PN0P_  (.D(_01780_),
    .DE(net299),
    .Q(\w[39][19] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][1]$_SDFFCE_PN0P_  (.D(_01781_),
    .DE(net298),
    .Q(\w[39][1] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][20]$_SDFFCE_PN0P_  (.D(_01782_),
    .DE(_00080_),
    .Q(\w[39][20] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][21]$_SDFFCE_PN0P_  (.D(_01783_),
    .DE(net299),
    .Q(\w[39][21] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][22]$_SDFFCE_PN0P_  (.D(_01784_),
    .DE(net299),
    .Q(\w[39][22] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][23]$_SDFFCE_PN0P_  (.D(_01785_),
    .DE(net300),
    .Q(\w[39][23] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][24]$_SDFFCE_PN0P_  (.D(_01786_),
    .DE(net300),
    .Q(\w[39][24] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][25]$_SDFFCE_PN0P_  (.D(_01787_),
    .DE(net299),
    .Q(\w[39][25] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][26]$_SDFFCE_PN0P_  (.D(_01788_),
    .DE(net298),
    .Q(\w[39][26] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][27]$_SDFFCE_PN0P_  (.D(_01789_),
    .DE(net300),
    .Q(\w[39][27] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][28]$_SDFFCE_PN0P_  (.D(_01790_),
    .DE(net298),
    .Q(\w[39][28] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][29]$_SDFFCE_PN0P_  (.D(_01791_),
    .DE(net300),
    .Q(\w[39][29] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][2]$_SDFFCE_PN0P_  (.D(_01792_),
    .DE(net298),
    .Q(\w[39][2] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][30]$_SDFFCE_PN0P_  (.D(_01793_),
    .DE(_00080_),
    .Q(\w[39][30] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][31]$_SDFFCE_PN0P_  (.D(_01794_),
    .DE(net298),
    .Q(\w[39][31] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][3]$_SDFFCE_PN0P_  (.D(_01795_),
    .DE(net298),
    .Q(\w[39][3] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][4]$_SDFFCE_PN0P_  (.D(_01796_),
    .DE(net300),
    .Q(\w[39][4] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][5]$_SDFFCE_PN0P_  (.D(_01797_),
    .DE(net298),
    .Q(\w[39][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][6]$_SDFFCE_PN0P_  (.D(_01798_),
    .DE(net299),
    .Q(\w[39][6] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][7]$_SDFFCE_PN0P_  (.D(_01799_),
    .DE(net298),
    .Q(\w[39][7] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][8]$_SDFFCE_PN0P_  (.D(_01800_),
    .DE(net300),
    .Q(\w[39][8] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[39][9]$_SDFFCE_PN0P_  (.D(_01801_),
    .DE(net300),
    .Q(\w[39][9] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][0]$_DFFE_PP_  (.D(_00417_),
    .DE(_00079_),
    .Q(\w[3][0] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][10]$_DFFE_PP_  (.D(_00418_),
    .DE(_00079_),
    .Q(\w[3][10] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][11]$_DFFE_PP_  (.D(_00419_),
    .DE(_00079_),
    .Q(\w[3][11] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][12]$_DFFE_PP_  (.D(_00420_),
    .DE(_00079_),
    .Q(\w[3][12] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][13]$_DFFE_PP_  (.D(_00421_),
    .DE(_00079_),
    .Q(\w[3][13] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][14]$_DFFE_PP_  (.D(_00422_),
    .DE(_00079_),
    .Q(\w[3][14] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][15]$_DFFE_PP_  (.D(_00423_),
    .DE(_00079_),
    .Q(\w[3][15] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][16]$_DFFE_PP_  (.D(_00424_),
    .DE(_00079_),
    .Q(\w[3][16] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][17]$_DFFE_PP_  (.D(_00425_),
    .DE(_00079_),
    .Q(\w[3][17] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][18]$_DFFE_PP_  (.D(_00426_),
    .DE(_00079_),
    .Q(\w[3][18] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][19]$_DFFE_PP_  (.D(_00427_),
    .DE(_00079_),
    .Q(\w[3][19] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][1]$_DFFE_PP_  (.D(_00428_),
    .DE(_00079_),
    .Q(\w[3][1] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][20]$_DFFE_PP_  (.D(_00429_),
    .DE(_00079_),
    .Q(\w[3][20] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][21]$_DFFE_PP_  (.D(_00430_),
    .DE(_00079_),
    .Q(\w[3][21] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][22]$_DFFE_PP_  (.D(_00431_),
    .DE(_00079_),
    .Q(\w[3][22] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][23]$_DFFE_PP_  (.D(_00432_),
    .DE(_00079_),
    .Q(\w[3][23] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][24]$_DFFE_PP_  (.D(_00433_),
    .DE(_00079_),
    .Q(\w[3][24] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][25]$_DFFE_PP_  (.D(_00434_),
    .DE(_00079_),
    .Q(\w[3][25] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][26]$_DFFE_PP_  (.D(_00435_),
    .DE(_00079_),
    .Q(\w[3][26] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][27]$_DFFE_PP_  (.D(_00436_),
    .DE(_00079_),
    .Q(\w[3][27] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][28]$_DFFE_PP_  (.D(_00437_),
    .DE(_00079_),
    .Q(\w[3][28] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][29]$_DFFE_PP_  (.D(_00438_),
    .DE(_00079_),
    .Q(\w[3][29] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][2]$_DFFE_PP_  (.D(_00439_),
    .DE(_00079_),
    .Q(\w[3][2] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][30]$_DFFE_PP_  (.D(_00440_),
    .DE(_00079_),
    .Q(\w[3][30] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][31]$_DFFE_PP_  (.D(_00441_),
    .DE(_00079_),
    .Q(\w[3][31] ),
    .CLK(clknet_leaf_289_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][3]$_DFFE_PP_  (.D(_00442_),
    .DE(_00079_),
    .Q(\w[3][3] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][4]$_DFFE_PP_  (.D(_00443_),
    .DE(_00079_),
    .Q(\w[3][4] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][5]$_DFFE_PP_  (.D(_00444_),
    .DE(_00079_),
    .Q(\w[3][5] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][6]$_DFFE_PP_  (.D(_00445_),
    .DE(_00079_),
    .Q(\w[3][6] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][7]$_DFFE_PP_  (.D(_00446_),
    .DE(_00079_),
    .Q(\w[3][7] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][8]$_DFFE_PP_  (.D(_00447_),
    .DE(_00079_),
    .Q(\w[3][8] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[3][9]$_DFFE_PP_  (.D(_00448_),
    .DE(_00079_),
    .Q(\w[3][9] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][0]$_SDFFCE_PN0P_  (.D(_01802_),
    .DE(_00110_),
    .Q(\w[40][0] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][10]$_SDFFCE_PN0P_  (.D(_01803_),
    .DE(_00110_),
    .Q(\w[40][10] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][11]$_SDFFCE_PN0P_  (.D(_01804_),
    .DE(_00110_),
    .Q(\w[40][11] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][12]$_SDFFCE_PN0P_  (.D(_01805_),
    .DE(_00110_),
    .Q(\w[40][12] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][13]$_SDFFCE_PN0P_  (.D(_01806_),
    .DE(_00110_),
    .Q(\w[40][13] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][14]$_SDFFCE_PN0P_  (.D(_01807_),
    .DE(_00110_),
    .Q(\w[40][14] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][15]$_SDFFCE_PN0P_  (.D(_01808_),
    .DE(_00110_),
    .Q(\w[40][15] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][16]$_SDFFCE_PN0P_  (.D(_01809_),
    .DE(_00110_),
    .Q(\w[40][16] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][17]$_SDFFCE_PN0P_  (.D(_01810_),
    .DE(_00110_),
    .Q(\w[40][17] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][18]$_SDFFCE_PN0P_  (.D(_01811_),
    .DE(_00110_),
    .Q(\w[40][18] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][19]$_SDFFCE_PN0P_  (.D(_01812_),
    .DE(_00110_),
    .Q(\w[40][19] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][1]$_SDFFCE_PN0P_  (.D(_01813_),
    .DE(_00110_),
    .Q(\w[40][1] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][20]$_SDFFCE_PN0P_  (.D(_01814_),
    .DE(_00110_),
    .Q(\w[40][20] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][21]$_SDFFCE_PN0P_  (.D(_01815_),
    .DE(_00110_),
    .Q(\w[40][21] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][22]$_SDFFCE_PN0P_  (.D(_01816_),
    .DE(_00110_),
    .Q(\w[40][22] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][23]$_SDFFCE_PN0P_  (.D(_01817_),
    .DE(_00110_),
    .Q(\w[40][23] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][24]$_SDFFCE_PN0P_  (.D(_01818_),
    .DE(_00110_),
    .Q(\w[40][24] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][25]$_SDFFCE_PN0P_  (.D(_01819_),
    .DE(_00110_),
    .Q(\w[40][25] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][26]$_SDFFCE_PN0P_  (.D(_01820_),
    .DE(_00110_),
    .Q(\w[40][26] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][27]$_SDFFCE_PN0P_  (.D(_01821_),
    .DE(_00110_),
    .Q(\w[40][27] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][28]$_SDFFCE_PN0P_  (.D(_01822_),
    .DE(_00110_),
    .Q(\w[40][28] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][29]$_SDFFCE_PN0P_  (.D(_01823_),
    .DE(_00110_),
    .Q(\w[40][29] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][2]$_SDFFCE_PN0P_  (.D(_01824_),
    .DE(_00110_),
    .Q(\w[40][2] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][30]$_SDFFCE_PN0P_  (.D(_01825_),
    .DE(_00110_),
    .Q(\w[40][30] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][31]$_SDFFCE_PN0P_  (.D(_01826_),
    .DE(_00110_),
    .Q(\w[40][31] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][3]$_SDFFCE_PN0P_  (.D(_01827_),
    .DE(_00110_),
    .Q(\w[40][3] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][4]$_SDFFCE_PN0P_  (.D(_01828_),
    .DE(_00110_),
    .Q(\w[40][4] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][5]$_SDFFCE_PN0P_  (.D(_01829_),
    .DE(_00110_),
    .Q(\w[40][5] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][6]$_SDFFCE_PN0P_  (.D(_01830_),
    .DE(_00110_),
    .Q(\w[40][6] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][7]$_SDFFCE_PN0P_  (.D(_01831_),
    .DE(_00110_),
    .Q(\w[40][7] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][8]$_SDFFCE_PN0P_  (.D(_01832_),
    .DE(_00110_),
    .Q(\w[40][8] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[40][9]$_SDFFCE_PN0P_  (.D(_01833_),
    .DE(_00110_),
    .Q(\w[40][9] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][0]$_SDFFCE_PN0P_  (.D(_01834_),
    .DE(_00078_),
    .Q(\w[41][0] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][10]$_SDFFCE_PN0P_  (.D(_01835_),
    .DE(_00078_),
    .Q(\w[41][10] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][11]$_SDFFCE_PN0P_  (.D(_01836_),
    .DE(_00078_),
    .Q(\w[41][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][12]$_SDFFCE_PN0P_  (.D(_01837_),
    .DE(_00078_),
    .Q(\w[41][12] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][13]$_SDFFCE_PN0P_  (.D(_01838_),
    .DE(_00078_),
    .Q(\w[41][13] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][14]$_SDFFCE_PN0P_  (.D(_01839_),
    .DE(_00078_),
    .Q(\w[41][14] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][15]$_SDFFCE_PN0P_  (.D(_01840_),
    .DE(_00078_),
    .Q(\w[41][15] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][16]$_SDFFCE_PN0P_  (.D(_01841_),
    .DE(_00078_),
    .Q(\w[41][16] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][17]$_SDFFCE_PN0P_  (.D(_01842_),
    .DE(_00078_),
    .Q(\w[41][17] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][18]$_SDFFCE_PN0P_  (.D(_01843_),
    .DE(_00078_),
    .Q(\w[41][18] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][19]$_SDFFCE_PN0P_  (.D(_01844_),
    .DE(_00078_),
    .Q(\w[41][19] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][1]$_SDFFCE_PN0P_  (.D(_01845_),
    .DE(_00078_),
    .Q(\w[41][1] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][20]$_SDFFCE_PN0P_  (.D(_01846_),
    .DE(_00078_),
    .Q(\w[41][20] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][21]$_SDFFCE_PN0P_  (.D(_01847_),
    .DE(_00078_),
    .Q(\w[41][21] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][22]$_SDFFCE_PN0P_  (.D(_01848_),
    .DE(_00078_),
    .Q(\w[41][22] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][23]$_SDFFCE_PN0P_  (.D(_01849_),
    .DE(_00078_),
    .Q(\w[41][23] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][24]$_SDFFCE_PN0P_  (.D(_01850_),
    .DE(_00078_),
    .Q(\w[41][24] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][25]$_SDFFCE_PN0P_  (.D(_01851_),
    .DE(_00078_),
    .Q(\w[41][25] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][26]$_SDFFCE_PN0P_  (.D(_01852_),
    .DE(_00078_),
    .Q(\w[41][26] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][27]$_SDFFCE_PN0P_  (.D(_01853_),
    .DE(_00078_),
    .Q(\w[41][27] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][28]$_SDFFCE_PN0P_  (.D(_01854_),
    .DE(_00078_),
    .Q(\w[41][28] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][29]$_SDFFCE_PN0P_  (.D(_01855_),
    .DE(_00078_),
    .Q(\w[41][29] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][2]$_SDFFCE_PN0P_  (.D(_01856_),
    .DE(_00078_),
    .Q(\w[41][2] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][30]$_SDFFCE_PN0P_  (.D(_01857_),
    .DE(_00078_),
    .Q(\w[41][30] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][31]$_SDFFCE_PN0P_  (.D(_01858_),
    .DE(_00078_),
    .Q(\w[41][31] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][3]$_SDFFCE_PN0P_  (.D(_01859_),
    .DE(_00078_),
    .Q(\w[41][3] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][4]$_SDFFCE_PN0P_  (.D(_01860_),
    .DE(_00078_),
    .Q(\w[41][4] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][5]$_SDFFCE_PN0P_  (.D(_01861_),
    .DE(_00078_),
    .Q(\w[41][5] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][6]$_SDFFCE_PN0P_  (.D(_01862_),
    .DE(_00078_),
    .Q(\w[41][6] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][7]$_SDFFCE_PN0P_  (.D(_01863_),
    .DE(_00078_),
    .Q(\w[41][7] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][8]$_SDFFCE_PN0P_  (.D(_01864_),
    .DE(_00078_),
    .Q(\w[41][8] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[41][9]$_SDFFCE_PN0P_  (.D(_01865_),
    .DE(_00078_),
    .Q(\w[41][9] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][0]$_SDFFCE_PN0P_  (.D(_01866_),
    .DE(_00109_),
    .Q(\w[42][0] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][10]$_SDFFCE_PN0P_  (.D(_01867_),
    .DE(_00109_),
    .Q(\w[42][10] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][11]$_SDFFCE_PN0P_  (.D(_01868_),
    .DE(_00109_),
    .Q(\w[42][11] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][12]$_SDFFCE_PN0P_  (.D(_01869_),
    .DE(_00109_),
    .Q(\w[42][12] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][13]$_SDFFCE_PN0P_  (.D(_01870_),
    .DE(_00109_),
    .Q(\w[42][13] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][14]$_SDFFCE_PN0P_  (.D(_01871_),
    .DE(_00109_),
    .Q(\w[42][14] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][15]$_SDFFCE_PN0P_  (.D(_01872_),
    .DE(_00109_),
    .Q(\w[42][15] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][16]$_SDFFCE_PN0P_  (.D(_01873_),
    .DE(_00109_),
    .Q(\w[42][16] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][17]$_SDFFCE_PN0P_  (.D(_01874_),
    .DE(_00109_),
    .Q(\w[42][17] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][18]$_SDFFCE_PN0P_  (.D(_01875_),
    .DE(_00109_),
    .Q(\w[42][18] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][19]$_SDFFCE_PN0P_  (.D(_01876_),
    .DE(_00109_),
    .Q(\w[42][19] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][1]$_SDFFCE_PN0P_  (.D(_01877_),
    .DE(_00109_),
    .Q(\w[42][1] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][20]$_SDFFCE_PN0P_  (.D(_01878_),
    .DE(_00109_),
    .Q(\w[42][20] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][21]$_SDFFCE_PN0P_  (.D(_01879_),
    .DE(_00109_),
    .Q(\w[42][21] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][22]$_SDFFCE_PN0P_  (.D(_01880_),
    .DE(_00109_),
    .Q(\w[42][22] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][23]$_SDFFCE_PN0P_  (.D(_01881_),
    .DE(_00109_),
    .Q(\w[42][23] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][24]$_SDFFCE_PN0P_  (.D(_01882_),
    .DE(_00109_),
    .Q(\w[42][24] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][25]$_SDFFCE_PN0P_  (.D(_01883_),
    .DE(_00109_),
    .Q(\w[42][25] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][26]$_SDFFCE_PN0P_  (.D(_01884_),
    .DE(_00109_),
    .Q(\w[42][26] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][27]$_SDFFCE_PN0P_  (.D(_01885_),
    .DE(_00109_),
    .Q(\w[42][27] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][28]$_SDFFCE_PN0P_  (.D(_01886_),
    .DE(_00109_),
    .Q(\w[42][28] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][29]$_SDFFCE_PN0P_  (.D(_01887_),
    .DE(_00109_),
    .Q(\w[42][29] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][2]$_SDFFCE_PN0P_  (.D(_01888_),
    .DE(_00109_),
    .Q(\w[42][2] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][30]$_SDFFCE_PN0P_  (.D(_01889_),
    .DE(_00109_),
    .Q(\w[42][30] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][31]$_SDFFCE_PN0P_  (.D(_01890_),
    .DE(_00109_),
    .Q(\w[42][31] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][3]$_SDFFCE_PN0P_  (.D(_01891_),
    .DE(_00109_),
    .Q(\w[42][3] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][4]$_SDFFCE_PN0P_  (.D(_01892_),
    .DE(_00109_),
    .Q(\w[42][4] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][5]$_SDFFCE_PN0P_  (.D(_01893_),
    .DE(_00109_),
    .Q(\w[42][5] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][6]$_SDFFCE_PN0P_  (.D(_01894_),
    .DE(_00109_),
    .Q(\w[42][6] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][7]$_SDFFCE_PN0P_  (.D(_01895_),
    .DE(_00109_),
    .Q(\w[42][7] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][8]$_SDFFCE_PN0P_  (.D(_01896_),
    .DE(_00109_),
    .Q(\w[42][8] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[42][9]$_SDFFCE_PN0P_  (.D(_01897_),
    .DE(_00109_),
    .Q(\w[42][9] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][0]$_SDFFCE_PN0P_  (.D(_01898_),
    .DE(_00077_),
    .Q(\w[43][0] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][10]$_SDFFCE_PN0P_  (.D(_01899_),
    .DE(_00077_),
    .Q(\w[43][10] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][11]$_SDFFCE_PN0P_  (.D(_01900_),
    .DE(_00077_),
    .Q(\w[43][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][12]$_SDFFCE_PN0P_  (.D(_01901_),
    .DE(_00077_),
    .Q(\w[43][12] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][13]$_SDFFCE_PN0P_  (.D(_01902_),
    .DE(_00077_),
    .Q(\w[43][13] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][14]$_SDFFCE_PN0P_  (.D(_01903_),
    .DE(_00077_),
    .Q(\w[43][14] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][15]$_SDFFCE_PN0P_  (.D(_01904_),
    .DE(_00077_),
    .Q(\w[43][15] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][16]$_SDFFCE_PN0P_  (.D(_01905_),
    .DE(_00077_),
    .Q(\w[43][16] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][17]$_SDFFCE_PN0P_  (.D(_01906_),
    .DE(_00077_),
    .Q(\w[43][17] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][18]$_SDFFCE_PN0P_  (.D(_01907_),
    .DE(_00077_),
    .Q(\w[43][18] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][19]$_SDFFCE_PN0P_  (.D(_01908_),
    .DE(_00077_),
    .Q(\w[43][19] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][1]$_SDFFCE_PN0P_  (.D(_01909_),
    .DE(_00077_),
    .Q(\w[43][1] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][20]$_SDFFCE_PN0P_  (.D(_01910_),
    .DE(_00077_),
    .Q(\w[43][20] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][21]$_SDFFCE_PN0P_  (.D(_01911_),
    .DE(_00077_),
    .Q(\w[43][21] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][22]$_SDFFCE_PN0P_  (.D(_01912_),
    .DE(_00077_),
    .Q(\w[43][22] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][23]$_SDFFCE_PN0P_  (.D(_01913_),
    .DE(_00077_),
    .Q(\w[43][23] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][24]$_SDFFCE_PN0P_  (.D(_01914_),
    .DE(_00077_),
    .Q(\w[43][24] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][25]$_SDFFCE_PN0P_  (.D(_01915_),
    .DE(_00077_),
    .Q(\w[43][25] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][26]$_SDFFCE_PN0P_  (.D(_01916_),
    .DE(_00077_),
    .Q(\w[43][26] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][27]$_SDFFCE_PN0P_  (.D(_01917_),
    .DE(_00077_),
    .Q(\w[43][27] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][28]$_SDFFCE_PN0P_  (.D(_01918_),
    .DE(_00077_),
    .Q(\w[43][28] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][29]$_SDFFCE_PN0P_  (.D(_01919_),
    .DE(_00077_),
    .Q(\w[43][29] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][2]$_SDFFCE_PN0P_  (.D(_01920_),
    .DE(_00077_),
    .Q(\w[43][2] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][30]$_SDFFCE_PN0P_  (.D(_01921_),
    .DE(_00077_),
    .Q(\w[43][30] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][31]$_SDFFCE_PN0P_  (.D(_01922_),
    .DE(_00077_),
    .Q(\w[43][31] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][3]$_SDFFCE_PN0P_  (.D(_01923_),
    .DE(_00077_),
    .Q(\w[43][3] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][4]$_SDFFCE_PN0P_  (.D(_01924_),
    .DE(_00077_),
    .Q(\w[43][4] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][5]$_SDFFCE_PN0P_  (.D(_01925_),
    .DE(_00077_),
    .Q(\w[43][5] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][6]$_SDFFCE_PN0P_  (.D(_01926_),
    .DE(_00077_),
    .Q(\w[43][6] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][7]$_SDFFCE_PN0P_  (.D(_01927_),
    .DE(_00077_),
    .Q(\w[43][7] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][8]$_SDFFCE_PN0P_  (.D(_01928_),
    .DE(_00077_),
    .Q(\w[43][8] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[43][9]$_SDFFCE_PN0P_  (.D(_01929_),
    .DE(_00077_),
    .Q(\w[43][9] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][0]$_SDFFCE_PN0P_  (.D(_01930_),
    .DE(_00108_),
    .Q(\w[44][0] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][10]$_SDFFCE_PN0P_  (.D(_01931_),
    .DE(_00108_),
    .Q(\w[44][10] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][11]$_SDFFCE_PN0P_  (.D(_01932_),
    .DE(_00108_),
    .Q(\w[44][11] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][12]$_SDFFCE_PN0P_  (.D(_01933_),
    .DE(_00108_),
    .Q(\w[44][12] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][13]$_SDFFCE_PN0P_  (.D(_01934_),
    .DE(_00108_),
    .Q(\w[44][13] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][14]$_SDFFCE_PN0P_  (.D(_01935_),
    .DE(_00108_),
    .Q(\w[44][14] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][15]$_SDFFCE_PN0P_  (.D(_01936_),
    .DE(_00108_),
    .Q(\w[44][15] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][16]$_SDFFCE_PN0P_  (.D(_01937_),
    .DE(_00108_),
    .Q(\w[44][16] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][17]$_SDFFCE_PN0P_  (.D(_01938_),
    .DE(_00108_),
    .Q(\w[44][17] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][18]$_SDFFCE_PN0P_  (.D(_01939_),
    .DE(_00108_),
    .Q(\w[44][18] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][19]$_SDFFCE_PN0P_  (.D(_01940_),
    .DE(_00108_),
    .Q(\w[44][19] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][1]$_SDFFCE_PN0P_  (.D(_01941_),
    .DE(_00108_),
    .Q(\w[44][1] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][20]$_SDFFCE_PN0P_  (.D(_01942_),
    .DE(_00108_),
    .Q(\w[44][20] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][21]$_SDFFCE_PN0P_  (.D(_01943_),
    .DE(_00108_),
    .Q(\w[44][21] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][22]$_SDFFCE_PN0P_  (.D(_01944_),
    .DE(_00108_),
    .Q(\w[44][22] ),
    .CLK(clknet_leaf_142_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][23]$_SDFFCE_PN0P_  (.D(_01945_),
    .DE(_00108_),
    .Q(\w[44][23] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][24]$_SDFFCE_PN0P_  (.D(_01946_),
    .DE(_00108_),
    .Q(\w[44][24] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][25]$_SDFFCE_PN0P_  (.D(_01947_),
    .DE(_00108_),
    .Q(\w[44][25] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][26]$_SDFFCE_PN0P_  (.D(_01948_),
    .DE(_00108_),
    .Q(\w[44][26] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][27]$_SDFFCE_PN0P_  (.D(_01949_),
    .DE(_00108_),
    .Q(\w[44][27] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][28]$_SDFFCE_PN0P_  (.D(_01950_),
    .DE(_00108_),
    .Q(\w[44][28] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][29]$_SDFFCE_PN0P_  (.D(_01951_),
    .DE(_00108_),
    .Q(\w[44][29] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][2]$_SDFFCE_PN0P_  (.D(_01952_),
    .DE(_00108_),
    .Q(\w[44][2] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][30]$_SDFFCE_PN0P_  (.D(_01953_),
    .DE(_00108_),
    .Q(\w[44][30] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][31]$_SDFFCE_PN0P_  (.D(_01954_),
    .DE(_00108_),
    .Q(\w[44][31] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][3]$_SDFFCE_PN0P_  (.D(_01955_),
    .DE(_00108_),
    .Q(\w[44][3] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][4]$_SDFFCE_PN0P_  (.D(_01956_),
    .DE(_00108_),
    .Q(\w[44][4] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][5]$_SDFFCE_PN0P_  (.D(_01957_),
    .DE(_00108_),
    .Q(\w[44][5] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][6]$_SDFFCE_PN0P_  (.D(_01958_),
    .DE(_00108_),
    .Q(\w[44][6] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][7]$_SDFFCE_PN0P_  (.D(_01959_),
    .DE(_00108_),
    .Q(\w[44][7] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][8]$_SDFFCE_PN0P_  (.D(_01960_),
    .DE(_00108_),
    .Q(\w[44][8] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[44][9]$_SDFFCE_PN0P_  (.D(_01961_),
    .DE(_00108_),
    .Q(\w[44][9] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][0]$_SDFFCE_PN0P_  (.D(_01962_),
    .DE(_00076_),
    .Q(\w[45][0] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][10]$_SDFFCE_PN0P_  (.D(_01963_),
    .DE(_00076_),
    .Q(\w[45][10] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][11]$_SDFFCE_PN0P_  (.D(_01964_),
    .DE(_00076_),
    .Q(\w[45][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][12]$_SDFFCE_PN0P_  (.D(_01965_),
    .DE(_00076_),
    .Q(\w[45][12] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][13]$_SDFFCE_PN0P_  (.D(_01966_),
    .DE(_00076_),
    .Q(\w[45][13] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][14]$_SDFFCE_PN0P_  (.D(_01967_),
    .DE(_00076_),
    .Q(\w[45][14] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][15]$_SDFFCE_PN0P_  (.D(_01968_),
    .DE(_00076_),
    .Q(\w[45][15] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][16]$_SDFFCE_PN0P_  (.D(_01969_),
    .DE(_00076_),
    .Q(\w[45][16] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][17]$_SDFFCE_PN0P_  (.D(_01970_),
    .DE(_00076_),
    .Q(\w[45][17] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][18]$_SDFFCE_PN0P_  (.D(_01971_),
    .DE(_00076_),
    .Q(\w[45][18] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][19]$_SDFFCE_PN0P_  (.D(_01972_),
    .DE(_00076_),
    .Q(\w[45][19] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][1]$_SDFFCE_PN0P_  (.D(_01973_),
    .DE(_00076_),
    .Q(\w[45][1] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][20]$_SDFFCE_PN0P_  (.D(_01974_),
    .DE(_00076_),
    .Q(\w[45][20] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][21]$_SDFFCE_PN0P_  (.D(_01975_),
    .DE(_00076_),
    .Q(\w[45][21] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][22]$_SDFFCE_PN0P_  (.D(_01976_),
    .DE(_00076_),
    .Q(\w[45][22] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][23]$_SDFFCE_PN0P_  (.D(_01977_),
    .DE(_00076_),
    .Q(\w[45][23] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][24]$_SDFFCE_PN0P_  (.D(_01978_),
    .DE(_00076_),
    .Q(\w[45][24] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][25]$_SDFFCE_PN0P_  (.D(_01979_),
    .DE(_00076_),
    .Q(\w[45][25] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][26]$_SDFFCE_PN0P_  (.D(_01980_),
    .DE(_00076_),
    .Q(\w[45][26] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][27]$_SDFFCE_PN0P_  (.D(_01981_),
    .DE(_00076_),
    .Q(\w[45][27] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][28]$_SDFFCE_PN0P_  (.D(_01982_),
    .DE(_00076_),
    .Q(\w[45][28] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][29]$_SDFFCE_PN0P_  (.D(_01983_),
    .DE(_00076_),
    .Q(\w[45][29] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][2]$_SDFFCE_PN0P_  (.D(_01984_),
    .DE(_00076_),
    .Q(\w[45][2] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][30]$_SDFFCE_PN0P_  (.D(_01985_),
    .DE(_00076_),
    .Q(\w[45][30] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][31]$_SDFFCE_PN0P_  (.D(_01986_),
    .DE(_00076_),
    .Q(\w[45][31] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][3]$_SDFFCE_PN0P_  (.D(_01987_),
    .DE(_00076_),
    .Q(\w[45][3] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][4]$_SDFFCE_PN0P_  (.D(_01988_),
    .DE(_00076_),
    .Q(\w[45][4] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][5]$_SDFFCE_PN0P_  (.D(_01989_),
    .DE(_00076_),
    .Q(\w[45][5] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][6]$_SDFFCE_PN0P_  (.D(_01990_),
    .DE(_00076_),
    .Q(\w[45][6] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][7]$_SDFFCE_PN0P_  (.D(_01991_),
    .DE(_00076_),
    .Q(\w[45][7] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][8]$_SDFFCE_PN0P_  (.D(_01992_),
    .DE(_00076_),
    .Q(\w[45][8] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[45][9]$_SDFFCE_PN0P_  (.D(_01993_),
    .DE(_00076_),
    .Q(\w[45][9] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][0]$_SDFFCE_PN0P_  (.D(_01994_),
    .DE(_00107_),
    .Q(\w[46][0] ),
    .CLK(clknet_leaf_129_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][10]$_SDFFCE_PN0P_  (.D(_01995_),
    .DE(_00107_),
    .Q(\w[46][10] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][11]$_SDFFCE_PN0P_  (.D(_01996_),
    .DE(_00107_),
    .Q(\w[46][11] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][12]$_SDFFCE_PN0P_  (.D(_01997_),
    .DE(_00107_),
    .Q(\w[46][12] ),
    .CLK(clknet_leaf_46_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][13]$_SDFFCE_PN0P_  (.D(_01998_),
    .DE(_00107_),
    .Q(\w[46][13] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][14]$_SDFFCE_PN0P_  (.D(_01999_),
    .DE(_00107_),
    .Q(\w[46][14] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][15]$_SDFFCE_PN0P_  (.D(_02000_),
    .DE(_00107_),
    .Q(\w[46][15] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][16]$_SDFFCE_PN0P_  (.D(_02001_),
    .DE(_00107_),
    .Q(\w[46][16] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][17]$_SDFFCE_PN0P_  (.D(_02002_),
    .DE(_00107_),
    .Q(\w[46][17] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][18]$_SDFFCE_PN0P_  (.D(_02003_),
    .DE(_00107_),
    .Q(\w[46][18] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][19]$_SDFFCE_PN0P_  (.D(_02004_),
    .DE(_00107_),
    .Q(\w[46][19] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][1]$_SDFFCE_PN0P_  (.D(_02005_),
    .DE(_00107_),
    .Q(\w[46][1] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][20]$_SDFFCE_PN0P_  (.D(_02006_),
    .DE(_00107_),
    .Q(\w[46][20] ),
    .CLK(clknet_leaf_177_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][21]$_SDFFCE_PN0P_  (.D(_02007_),
    .DE(_00107_),
    .Q(\w[46][21] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][22]$_SDFFCE_PN0P_  (.D(_02008_),
    .DE(_00107_),
    .Q(\w[46][22] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][23]$_SDFFCE_PN0P_  (.D(_02009_),
    .DE(_00107_),
    .Q(\w[46][23] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][24]$_SDFFCE_PN0P_  (.D(_02010_),
    .DE(_00107_),
    .Q(\w[46][24] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][25]$_SDFFCE_PN0P_  (.D(_02011_),
    .DE(_00107_),
    .Q(\w[46][25] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][26]$_SDFFCE_PN0P_  (.D(_02012_),
    .DE(_00107_),
    .Q(\w[46][26] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][27]$_SDFFCE_PN0P_  (.D(_02013_),
    .DE(_00107_),
    .Q(\w[46][27] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][28]$_SDFFCE_PN0P_  (.D(_02014_),
    .DE(_00107_),
    .Q(\w[46][28] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][29]$_SDFFCE_PN0P_  (.D(_02015_),
    .DE(_00107_),
    .Q(\w[46][29] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][2]$_SDFFCE_PN0P_  (.D(_02016_),
    .DE(_00107_),
    .Q(\w[46][2] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][30]$_SDFFCE_PN0P_  (.D(_02017_),
    .DE(_00107_),
    .Q(\w[46][30] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][31]$_SDFFCE_PN0P_  (.D(_02018_),
    .DE(_00107_),
    .Q(\w[46][31] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][3]$_SDFFCE_PN0P_  (.D(_02019_),
    .DE(_00107_),
    .Q(\w[46][3] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][4]$_SDFFCE_PN0P_  (.D(_02020_),
    .DE(_00107_),
    .Q(\w[46][4] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][5]$_SDFFCE_PN0P_  (.D(_02021_),
    .DE(_00107_),
    .Q(\w[46][5] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][6]$_SDFFCE_PN0P_  (.D(_02022_),
    .DE(_00107_),
    .Q(\w[46][6] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][7]$_SDFFCE_PN0P_  (.D(_02023_),
    .DE(_00107_),
    .Q(\w[46][7] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][8]$_SDFFCE_PN0P_  (.D(_02024_),
    .DE(_00107_),
    .Q(\w[46][8] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[46][9]$_SDFFCE_PN0P_  (.D(_02025_),
    .DE(_00107_),
    .Q(\w[46][9] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][0]$_SDFFCE_PN0P_  (.D(_02026_),
    .DE(_00075_),
    .Q(\w[47][0] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][10]$_SDFFCE_PN0P_  (.D(_02027_),
    .DE(_00075_),
    .Q(\w[47][10] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][11]$_SDFFCE_PN0P_  (.D(_02028_),
    .DE(_00075_),
    .Q(\w[47][11] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][12]$_SDFFCE_PN0P_  (.D(_02029_),
    .DE(_00075_),
    .Q(\w[47][12] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][13]$_SDFFCE_PN0P_  (.D(_02030_),
    .DE(_00075_),
    .Q(\w[47][13] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][14]$_SDFFCE_PN0P_  (.D(_02031_),
    .DE(_00075_),
    .Q(\w[47][14] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][15]$_SDFFCE_PN0P_  (.D(_02032_),
    .DE(_00075_),
    .Q(\w[47][15] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][16]$_SDFFCE_PN0P_  (.D(_02033_),
    .DE(_00075_),
    .Q(\w[47][16] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][17]$_SDFFCE_PN0P_  (.D(_02034_),
    .DE(_00075_),
    .Q(\w[47][17] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][18]$_SDFFCE_PN0P_  (.D(_02035_),
    .DE(_00075_),
    .Q(\w[47][18] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][19]$_SDFFCE_PN0P_  (.D(_02036_),
    .DE(_00075_),
    .Q(\w[47][19] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][1]$_SDFFCE_PN0P_  (.D(_02037_),
    .DE(_00075_),
    .Q(\w[47][1] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][20]$_SDFFCE_PN0P_  (.D(_02038_),
    .DE(_00075_),
    .Q(\w[47][20] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][21]$_SDFFCE_PN0P_  (.D(_02039_),
    .DE(_00075_),
    .Q(\w[47][21] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][22]$_SDFFCE_PN0P_  (.D(_02040_),
    .DE(_00075_),
    .Q(\w[47][22] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][23]$_SDFFCE_PN0P_  (.D(_02041_),
    .DE(_00075_),
    .Q(\w[47][23] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][24]$_SDFFCE_PN0P_  (.D(_02042_),
    .DE(_00075_),
    .Q(\w[47][24] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][25]$_SDFFCE_PN0P_  (.D(_02043_),
    .DE(_00075_),
    .Q(\w[47][25] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][26]$_SDFFCE_PN0P_  (.D(_02044_),
    .DE(_00075_),
    .Q(\w[47][26] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][27]$_SDFFCE_PN0P_  (.D(_02045_),
    .DE(_00075_),
    .Q(\w[47][27] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][28]$_SDFFCE_PN0P_  (.D(_02046_),
    .DE(_00075_),
    .Q(\w[47][28] ),
    .CLK(clknet_leaf_15_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][29]$_SDFFCE_PN0P_  (.D(_02047_),
    .DE(_00075_),
    .Q(\w[47][29] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][2]$_SDFFCE_PN0P_  (.D(_02048_),
    .DE(_00075_),
    .Q(\w[47][2] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][30]$_SDFFCE_PN0P_  (.D(_02049_),
    .DE(_00075_),
    .Q(\w[47][30] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][31]$_SDFFCE_PN0P_  (.D(_02050_),
    .DE(_00075_),
    .Q(\w[47][31] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][3]$_SDFFCE_PN0P_  (.D(_02051_),
    .DE(_00075_),
    .Q(\w[47][3] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][4]$_SDFFCE_PN0P_  (.D(_02052_),
    .DE(_00075_),
    .Q(\w[47][4] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][5]$_SDFFCE_PN0P_  (.D(_02053_),
    .DE(_00075_),
    .Q(\w[47][5] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][6]$_SDFFCE_PN0P_  (.D(_02054_),
    .DE(_00075_),
    .Q(\w[47][6] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][7]$_SDFFCE_PN0P_  (.D(_02055_),
    .DE(_00075_),
    .Q(\w[47][7] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][8]$_SDFFCE_PN0P_  (.D(_02056_),
    .DE(_00075_),
    .Q(\w[47][8] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[47][9]$_SDFFCE_PN0P_  (.D(_02057_),
    .DE(_00075_),
    .Q(\w[47][9] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][0]$_SDFFCE_PN0P_  (.D(_02058_),
    .DE(_00106_),
    .Q(\w[48][0] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][10]$_SDFFCE_PN0P_  (.D(_02059_),
    .DE(_00106_),
    .Q(\w[48][10] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][11]$_SDFFCE_PN0P_  (.D(_02060_),
    .DE(_00106_),
    .Q(\w[48][11] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][12]$_SDFFCE_PN0P_  (.D(_02061_),
    .DE(_00106_),
    .Q(\w[48][12] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][13]$_SDFFCE_PN0P_  (.D(_02062_),
    .DE(_00106_),
    .Q(\w[48][13] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][14]$_SDFFCE_PN0P_  (.D(_02063_),
    .DE(_00106_),
    .Q(\w[48][14] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][15]$_SDFFCE_PN0P_  (.D(_02064_),
    .DE(_00106_),
    .Q(\w[48][15] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][16]$_SDFFCE_PN0P_  (.D(_02065_),
    .DE(_00106_),
    .Q(\w[48][16] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][17]$_SDFFCE_PN0P_  (.D(_02066_),
    .DE(_00106_),
    .Q(\w[48][17] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][18]$_SDFFCE_PN0P_  (.D(_02067_),
    .DE(_00106_),
    .Q(\w[48][18] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][19]$_SDFFCE_PN0P_  (.D(_02068_),
    .DE(_00106_),
    .Q(\w[48][19] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][1]$_SDFFCE_PN0P_  (.D(_02069_),
    .DE(_00106_),
    .Q(\w[48][1] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][20]$_SDFFCE_PN0P_  (.D(_02070_),
    .DE(_00106_),
    .Q(\w[48][20] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][21]$_SDFFCE_PN0P_  (.D(_02071_),
    .DE(_00106_),
    .Q(\w[48][21] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][22]$_SDFFCE_PN0P_  (.D(_02072_),
    .DE(_00106_),
    .Q(\w[48][22] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][23]$_SDFFCE_PN0P_  (.D(_02073_),
    .DE(_00106_),
    .Q(\w[48][23] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][24]$_SDFFCE_PN0P_  (.D(_02074_),
    .DE(_00106_),
    .Q(\w[48][24] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][25]$_SDFFCE_PN0P_  (.D(_02075_),
    .DE(_00106_),
    .Q(\w[48][25] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][26]$_SDFFCE_PN0P_  (.D(_02076_),
    .DE(_00106_),
    .Q(\w[48][26] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][27]$_SDFFCE_PN0P_  (.D(_02077_),
    .DE(_00106_),
    .Q(\w[48][27] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][28]$_SDFFCE_PN0P_  (.D(_02078_),
    .DE(_00106_),
    .Q(\w[48][28] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][29]$_SDFFCE_PN0P_  (.D(_02079_),
    .DE(_00106_),
    .Q(\w[48][29] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][2]$_SDFFCE_PN0P_  (.D(_02080_),
    .DE(_00106_),
    .Q(\w[48][2] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][30]$_SDFFCE_PN0P_  (.D(_02081_),
    .DE(_00106_),
    .Q(\w[48][30] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][31]$_SDFFCE_PN0P_  (.D(_02082_),
    .DE(_00106_),
    .Q(\w[48][31] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][3]$_SDFFCE_PN0P_  (.D(_02083_),
    .DE(_00106_),
    .Q(\w[48][3] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][4]$_SDFFCE_PN0P_  (.D(_02084_),
    .DE(_00106_),
    .Q(\w[48][4] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][5]$_SDFFCE_PN0P_  (.D(_02085_),
    .DE(_00106_),
    .Q(\w[48][5] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][6]$_SDFFCE_PN0P_  (.D(_02086_),
    .DE(_00106_),
    .Q(\w[48][6] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][7]$_SDFFCE_PN0P_  (.D(_02087_),
    .DE(_00106_),
    .Q(\w[48][7] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][8]$_SDFFCE_PN0P_  (.D(_02088_),
    .DE(_00106_),
    .Q(\w[48][8] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[48][9]$_SDFFCE_PN0P_  (.D(_02089_),
    .DE(_00106_),
    .Q(\w[48][9] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][0]$_SDFFCE_PN0P_  (.D(_02090_),
    .DE(_00074_),
    .Q(\w[49][0] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][10]$_SDFFCE_PN0P_  (.D(_02091_),
    .DE(_00074_),
    .Q(\w[49][10] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][11]$_SDFFCE_PN0P_  (.D(_02092_),
    .DE(_00074_),
    .Q(\w[49][11] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][12]$_SDFFCE_PN0P_  (.D(_02093_),
    .DE(_00074_),
    .Q(\w[49][12] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][13]$_SDFFCE_PN0P_  (.D(_02094_),
    .DE(_00074_),
    .Q(\w[49][13] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][14]$_SDFFCE_PN0P_  (.D(_02095_),
    .DE(_00074_),
    .Q(\w[49][14] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][15]$_SDFFCE_PN0P_  (.D(_02096_),
    .DE(_00074_),
    .Q(\w[49][15] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][16]$_SDFFCE_PN0P_  (.D(_02097_),
    .DE(_00074_),
    .Q(\w[49][16] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][17]$_SDFFCE_PN0P_  (.D(_02098_),
    .DE(_00074_),
    .Q(\w[49][17] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][18]$_SDFFCE_PN0P_  (.D(_02099_),
    .DE(_00074_),
    .Q(\w[49][18] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][19]$_SDFFCE_PN0P_  (.D(_02100_),
    .DE(_00074_),
    .Q(\w[49][19] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][1]$_SDFFCE_PN0P_  (.D(_02101_),
    .DE(_00074_),
    .Q(\w[49][1] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][20]$_SDFFCE_PN0P_  (.D(_02102_),
    .DE(_00074_),
    .Q(\w[49][20] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][21]$_SDFFCE_PN0P_  (.D(_02103_),
    .DE(_00074_),
    .Q(\w[49][21] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][22]$_SDFFCE_PN0P_  (.D(_02104_),
    .DE(_00074_),
    .Q(\w[49][22] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][23]$_SDFFCE_PN0P_  (.D(_02105_),
    .DE(_00074_),
    .Q(\w[49][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][24]$_SDFFCE_PN0P_  (.D(_02106_),
    .DE(_00074_),
    .Q(\w[49][24] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][25]$_SDFFCE_PN0P_  (.D(_02107_),
    .DE(_00074_),
    .Q(\w[49][25] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][26]$_SDFFCE_PN0P_  (.D(_02108_),
    .DE(_00074_),
    .Q(\w[49][26] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][27]$_SDFFCE_PN0P_  (.D(_02109_),
    .DE(_00074_),
    .Q(\w[49][27] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][28]$_SDFFCE_PN0P_  (.D(_02110_),
    .DE(_00074_),
    .Q(\w[49][28] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][29]$_SDFFCE_PN0P_  (.D(_02111_),
    .DE(_00074_),
    .Q(\w[49][29] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][2]$_SDFFCE_PN0P_  (.D(_02112_),
    .DE(_00074_),
    .Q(\w[49][2] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][30]$_SDFFCE_PN0P_  (.D(_02113_),
    .DE(_00074_),
    .Q(\w[49][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][31]$_SDFFCE_PN0P_  (.D(_02114_),
    .DE(_00074_),
    .Q(\w[49][31] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][3]$_SDFFCE_PN0P_  (.D(_02115_),
    .DE(_00074_),
    .Q(\w[49][3] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][4]$_SDFFCE_PN0P_  (.D(_02116_),
    .DE(_00074_),
    .Q(\w[49][4] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][5]$_SDFFCE_PN0P_  (.D(_02117_),
    .DE(_00074_),
    .Q(\w[49][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][6]$_SDFFCE_PN0P_  (.D(_02118_),
    .DE(_00074_),
    .Q(\w[49][6] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][7]$_SDFFCE_PN0P_  (.D(_02119_),
    .DE(_00074_),
    .Q(\w[49][7] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][8]$_SDFFCE_PN0P_  (.D(_02120_),
    .DE(_00074_),
    .Q(\w[49][8] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[49][9]$_SDFFCE_PN0P_  (.D(_02121_),
    .DE(_00074_),
    .Q(\w[49][9] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][0]$_DFFE_PP_  (.D(_00449_),
    .DE(_00105_),
    .Q(\w[4][0] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][10]$_DFFE_PP_  (.D(_00450_),
    .DE(_00105_),
    .Q(\w[4][10] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][11]$_DFFE_PP_  (.D(_00451_),
    .DE(_00105_),
    .Q(\w[4][11] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][12]$_DFFE_PP_  (.D(_00452_),
    .DE(_00105_),
    .Q(\w[4][12] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][13]$_DFFE_PP_  (.D(_00453_),
    .DE(_00105_),
    .Q(\w[4][13] ),
    .CLK(clknet_leaf_88_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][14]$_DFFE_PP_  (.D(_00454_),
    .DE(_00105_),
    .Q(\w[4][14] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][15]$_DFFE_PP_  (.D(_00455_),
    .DE(_00105_),
    .Q(\w[4][15] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][16]$_DFFE_PP_  (.D(_00456_),
    .DE(_00105_),
    .Q(\w[4][16] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][17]$_DFFE_PP_  (.D(_00457_),
    .DE(_00105_),
    .Q(\w[4][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][18]$_DFFE_PP_  (.D(_00458_),
    .DE(_00105_),
    .Q(\w[4][18] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][19]$_DFFE_PP_  (.D(_00459_),
    .DE(_00105_),
    .Q(\w[4][19] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][1]$_DFFE_PP_  (.D(_00460_),
    .DE(_00105_),
    .Q(\w[4][1] ),
    .CLK(clknet_leaf_143_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][20]$_DFFE_PP_  (.D(_00461_),
    .DE(_00105_),
    .Q(\w[4][20] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][21]$_DFFE_PP_  (.D(_00462_),
    .DE(_00105_),
    .Q(\w[4][21] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][22]$_DFFE_PP_  (.D(_00463_),
    .DE(_00105_),
    .Q(\w[4][22] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][23]$_DFFE_PP_  (.D(_00464_),
    .DE(_00105_),
    .Q(\w[4][23] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][24]$_DFFE_PP_  (.D(_00465_),
    .DE(_00105_),
    .Q(\w[4][24] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][25]$_DFFE_PP_  (.D(_00466_),
    .DE(_00105_),
    .Q(\w[4][25] ),
    .CLK(clknet_leaf_101_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][26]$_DFFE_PP_  (.D(_00467_),
    .DE(_00105_),
    .Q(\w[4][26] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][27]$_DFFE_PP_  (.D(_00468_),
    .DE(_00105_),
    .Q(\w[4][27] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][28]$_DFFE_PP_  (.D(_00469_),
    .DE(_00105_),
    .Q(\w[4][28] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][29]$_DFFE_PP_  (.D(_00470_),
    .DE(_00105_),
    .Q(\w[4][29] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][2]$_DFFE_PP_  (.D(_00471_),
    .DE(_00105_),
    .Q(\w[4][2] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][30]$_DFFE_PP_  (.D(_00472_),
    .DE(_00105_),
    .Q(\w[4][30] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][31]$_DFFE_PP_  (.D(_00473_),
    .DE(_00105_),
    .Q(\w[4][31] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][3]$_DFFE_PP_  (.D(_00474_),
    .DE(_00105_),
    .Q(\w[4][3] ),
    .CLK(clknet_leaf_56_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][4]$_DFFE_PP_  (.D(_00475_),
    .DE(_00105_),
    .Q(\w[4][4] ),
    .CLK(clknet_leaf_73_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][5]$_DFFE_PP_  (.D(_00476_),
    .DE(_00105_),
    .Q(\w[4][5] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][6]$_DFFE_PP_  (.D(_00477_),
    .DE(_00105_),
    .Q(\w[4][6] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][7]$_DFFE_PP_  (.D(_00478_),
    .DE(_00105_),
    .Q(\w[4][7] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][8]$_DFFE_PP_  (.D(_00479_),
    .DE(_00105_),
    .Q(\w[4][8] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[4][9]$_DFFE_PP_  (.D(_00480_),
    .DE(_00105_),
    .Q(\w[4][9] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][0]$_SDFFCE_PN0P_  (.D(_02122_),
    .DE(_00104_),
    .Q(\w[50][0] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][10]$_SDFFCE_PN0P_  (.D(_02123_),
    .DE(_00104_),
    .Q(\w[50][10] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][11]$_SDFFCE_PN0P_  (.D(_02124_),
    .DE(_00104_),
    .Q(\w[50][11] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][12]$_SDFFCE_PN0P_  (.D(_02125_),
    .DE(_00104_),
    .Q(\w[50][12] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][13]$_SDFFCE_PN0P_  (.D(_02126_),
    .DE(_00104_),
    .Q(\w[50][13] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][14]$_SDFFCE_PN0P_  (.D(_02127_),
    .DE(_00104_),
    .Q(\w[50][14] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][15]$_SDFFCE_PN0P_  (.D(_02128_),
    .DE(_00104_),
    .Q(\w[50][15] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][16]$_SDFFCE_PN0P_  (.D(_02129_),
    .DE(_00104_),
    .Q(\w[50][16] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][17]$_SDFFCE_PN0P_  (.D(_02130_),
    .DE(_00104_),
    .Q(\w[50][17] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][18]$_SDFFCE_PN0P_  (.D(_02131_),
    .DE(_00104_),
    .Q(\w[50][18] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][19]$_SDFFCE_PN0P_  (.D(_02132_),
    .DE(_00104_),
    .Q(\w[50][19] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][1]$_SDFFCE_PN0P_  (.D(_02133_),
    .DE(_00104_),
    .Q(\w[50][1] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][20]$_SDFFCE_PN0P_  (.D(_02134_),
    .DE(_00104_),
    .Q(\w[50][20] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][21]$_SDFFCE_PN0P_  (.D(_02135_),
    .DE(_00104_),
    .Q(\w[50][21] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][22]$_SDFFCE_PN0P_  (.D(_02136_),
    .DE(_00104_),
    .Q(\w[50][22] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][23]$_SDFFCE_PN0P_  (.D(_02137_),
    .DE(_00104_),
    .Q(\w[50][23] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][24]$_SDFFCE_PN0P_  (.D(_02138_),
    .DE(_00104_),
    .Q(\w[50][24] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][25]$_SDFFCE_PN0P_  (.D(_02139_),
    .DE(_00104_),
    .Q(\w[50][25] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][26]$_SDFFCE_PN0P_  (.D(_02140_),
    .DE(_00104_),
    .Q(\w[50][26] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][27]$_SDFFCE_PN0P_  (.D(_02141_),
    .DE(_00104_),
    .Q(\w[50][27] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][28]$_SDFFCE_PN0P_  (.D(_02142_),
    .DE(_00104_),
    .Q(\w[50][28] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][29]$_SDFFCE_PN0P_  (.D(_02143_),
    .DE(_00104_),
    .Q(\w[50][29] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][2]$_SDFFCE_PN0P_  (.D(_02144_),
    .DE(_00104_),
    .Q(\w[50][2] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][30]$_SDFFCE_PN0P_  (.D(_02145_),
    .DE(_00104_),
    .Q(\w[50][30] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][31]$_SDFFCE_PN0P_  (.D(_02146_),
    .DE(_00104_),
    .Q(\w[50][31] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][3]$_SDFFCE_PN0P_  (.D(_02147_),
    .DE(_00104_),
    .Q(\w[50][3] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][4]$_SDFFCE_PN0P_  (.D(_02148_),
    .DE(_00104_),
    .Q(\w[50][4] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][5]$_SDFFCE_PN0P_  (.D(_02149_),
    .DE(_00104_),
    .Q(\w[50][5] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][6]$_SDFFCE_PN0P_  (.D(_02150_),
    .DE(_00104_),
    .Q(\w[50][6] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][7]$_SDFFCE_PN0P_  (.D(_02151_),
    .DE(_00104_),
    .Q(\w[50][7] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][8]$_SDFFCE_PN0P_  (.D(_02152_),
    .DE(_00104_),
    .Q(\w[50][8] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[50][9]$_SDFFCE_PN0P_  (.D(_02153_),
    .DE(_00104_),
    .Q(\w[50][9] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][0]$_SDFFCE_PN0P_  (.D(_02154_),
    .DE(_00073_),
    .Q(\w[51][0] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][10]$_SDFFCE_PN0P_  (.D(_02155_),
    .DE(_00073_),
    .Q(\w[51][10] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][11]$_SDFFCE_PN0P_  (.D(_02156_),
    .DE(_00073_),
    .Q(\w[51][11] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][12]$_SDFFCE_PN0P_  (.D(_02157_),
    .DE(_00073_),
    .Q(\w[51][12] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][13]$_SDFFCE_PN0P_  (.D(_02158_),
    .DE(_00073_),
    .Q(\w[51][13] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][14]$_SDFFCE_PN0P_  (.D(_02159_),
    .DE(_00073_),
    .Q(\w[51][14] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][15]$_SDFFCE_PN0P_  (.D(_02160_),
    .DE(_00073_),
    .Q(\w[51][15] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][16]$_SDFFCE_PN0P_  (.D(_02161_),
    .DE(_00073_),
    .Q(\w[51][16] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][17]$_SDFFCE_PN0P_  (.D(_02162_),
    .DE(_00073_),
    .Q(\w[51][17] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][18]$_SDFFCE_PN0P_  (.D(_02163_),
    .DE(_00073_),
    .Q(\w[51][18] ),
    .CLK(clknet_leaf_229_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][19]$_SDFFCE_PN0P_  (.D(_02164_),
    .DE(_00073_),
    .Q(\w[51][19] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][1]$_SDFFCE_PN0P_  (.D(_02165_),
    .DE(_00073_),
    .Q(\w[51][1] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][20]$_SDFFCE_PN0P_  (.D(_02166_),
    .DE(_00073_),
    .Q(\w[51][20] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][21]$_SDFFCE_PN0P_  (.D(_02167_),
    .DE(_00073_),
    .Q(\w[51][21] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][22]$_SDFFCE_PN0P_  (.D(_02168_),
    .DE(_00073_),
    .Q(\w[51][22] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][23]$_SDFFCE_PN0P_  (.D(_02169_),
    .DE(_00073_),
    .Q(\w[51][23] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][24]$_SDFFCE_PN0P_  (.D(_02170_),
    .DE(_00073_),
    .Q(\w[51][24] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][25]$_SDFFCE_PN0P_  (.D(_02171_),
    .DE(_00073_),
    .Q(\w[51][25] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][26]$_SDFFCE_PN0P_  (.D(_02172_),
    .DE(_00073_),
    .Q(\w[51][26] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][27]$_SDFFCE_PN0P_  (.D(_02173_),
    .DE(_00073_),
    .Q(\w[51][27] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][28]$_SDFFCE_PN0P_  (.D(_02174_),
    .DE(_00073_),
    .Q(\w[51][28] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][29]$_SDFFCE_PN0P_  (.D(_02175_),
    .DE(_00073_),
    .Q(\w[51][29] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][2]$_SDFFCE_PN0P_  (.D(_02176_),
    .DE(_00073_),
    .Q(\w[51][2] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][30]$_SDFFCE_PN0P_  (.D(_02177_),
    .DE(_00073_),
    .Q(\w[51][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][31]$_SDFFCE_PN0P_  (.D(_02178_),
    .DE(_00073_),
    .Q(\w[51][31] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][3]$_SDFFCE_PN0P_  (.D(_02179_),
    .DE(_00073_),
    .Q(\w[51][3] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][4]$_SDFFCE_PN0P_  (.D(_02180_),
    .DE(_00073_),
    .Q(\w[51][4] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][5]$_SDFFCE_PN0P_  (.D(_02181_),
    .DE(_00073_),
    .Q(\w[51][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][6]$_SDFFCE_PN0P_  (.D(_02182_),
    .DE(_00073_),
    .Q(\w[51][6] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][7]$_SDFFCE_PN0P_  (.D(_02183_),
    .DE(_00073_),
    .Q(\w[51][7] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][8]$_SDFFCE_PN0P_  (.D(_02184_),
    .DE(_00073_),
    .Q(\w[51][8] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[51][9]$_SDFFCE_PN0P_  (.D(_02185_),
    .DE(_00073_),
    .Q(\w[51][9] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][0]$_SDFFCE_PN0P_  (.D(_02186_),
    .DE(_00103_),
    .Q(\w[52][0] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][10]$_SDFFCE_PN0P_  (.D(_02187_),
    .DE(_00103_),
    .Q(\w[52][10] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][11]$_SDFFCE_PN0P_  (.D(_02188_),
    .DE(_00103_),
    .Q(\w[52][11] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][12]$_SDFFCE_PN0P_  (.D(_02189_),
    .DE(_00103_),
    .Q(\w[52][12] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][13]$_SDFFCE_PN0P_  (.D(_02190_),
    .DE(_00103_),
    .Q(\w[52][13] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][14]$_SDFFCE_PN0P_  (.D(_02191_),
    .DE(_00103_),
    .Q(\w[52][14] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][15]$_SDFFCE_PN0P_  (.D(_02192_),
    .DE(_00103_),
    .Q(\w[52][15] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][16]$_SDFFCE_PN0P_  (.D(_02193_),
    .DE(_00103_),
    .Q(\w[52][16] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][17]$_SDFFCE_PN0P_  (.D(_02194_),
    .DE(_00103_),
    .Q(\w[52][17] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][18]$_SDFFCE_PN0P_  (.D(_02195_),
    .DE(_00103_),
    .Q(\w[52][18] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][19]$_SDFFCE_PN0P_  (.D(_02196_),
    .DE(_00103_),
    .Q(\w[52][19] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][1]$_SDFFCE_PN0P_  (.D(_02197_),
    .DE(_00103_),
    .Q(\w[52][1] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][20]$_SDFFCE_PN0P_  (.D(_02198_),
    .DE(_00103_),
    .Q(\w[52][20] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][21]$_SDFFCE_PN0P_  (.D(_02199_),
    .DE(_00103_),
    .Q(\w[52][21] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][22]$_SDFFCE_PN0P_  (.D(_02200_),
    .DE(_00103_),
    .Q(\w[52][22] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][23]$_SDFFCE_PN0P_  (.D(_02201_),
    .DE(_00103_),
    .Q(\w[52][23] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][24]$_SDFFCE_PN0P_  (.D(_02202_),
    .DE(_00103_),
    .Q(\w[52][24] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][25]$_SDFFCE_PN0P_  (.D(_02203_),
    .DE(_00103_),
    .Q(\w[52][25] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][26]$_SDFFCE_PN0P_  (.D(_02204_),
    .DE(_00103_),
    .Q(\w[52][26] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][27]$_SDFFCE_PN0P_  (.D(_02205_),
    .DE(_00103_),
    .Q(\w[52][27] ),
    .CLK(clknet_leaf_85_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][28]$_SDFFCE_PN0P_  (.D(_02206_),
    .DE(_00103_),
    .Q(\w[52][28] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][29]$_SDFFCE_PN0P_  (.D(_02207_),
    .DE(_00103_),
    .Q(\w[52][29] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][2]$_SDFFCE_PN0P_  (.D(_02208_),
    .DE(_00103_),
    .Q(\w[52][2] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][30]$_SDFFCE_PN0P_  (.D(_02209_),
    .DE(_00103_),
    .Q(\w[52][30] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][31]$_SDFFCE_PN0P_  (.D(_02210_),
    .DE(_00103_),
    .Q(\w[52][31] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][3]$_SDFFCE_PN0P_  (.D(_02211_),
    .DE(_00103_),
    .Q(\w[52][3] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][4]$_SDFFCE_PN0P_  (.D(_02212_),
    .DE(_00103_),
    .Q(\w[52][4] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][5]$_SDFFCE_PN0P_  (.D(_02213_),
    .DE(_00103_),
    .Q(\w[52][5] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][6]$_SDFFCE_PN0P_  (.D(_02214_),
    .DE(_00103_),
    .Q(\w[52][6] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][7]$_SDFFCE_PN0P_  (.D(_02215_),
    .DE(_00103_),
    .Q(\w[52][7] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][8]$_SDFFCE_PN0P_  (.D(_02216_),
    .DE(_00103_),
    .Q(\w[52][8] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[52][9]$_SDFFCE_PN0P_  (.D(_02217_),
    .DE(_00103_),
    .Q(\w[52][9] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][0]$_SDFFCE_PN0P_  (.D(_02218_),
    .DE(_00072_),
    .Q(\w[53][0] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][10]$_SDFFCE_PN0P_  (.D(_02219_),
    .DE(_00072_),
    .Q(\w[53][10] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][11]$_SDFFCE_PN0P_  (.D(_02220_),
    .DE(_00072_),
    .Q(\w[53][11] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][12]$_SDFFCE_PN0P_  (.D(_02221_),
    .DE(_00072_),
    .Q(\w[53][12] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][13]$_SDFFCE_PN0P_  (.D(_02222_),
    .DE(_00072_),
    .Q(\w[53][13] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][14]$_SDFFCE_PN0P_  (.D(_02223_),
    .DE(_00072_),
    .Q(\w[53][14] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][15]$_SDFFCE_PN0P_  (.D(_02224_),
    .DE(_00072_),
    .Q(\w[53][15] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][16]$_SDFFCE_PN0P_  (.D(_02225_),
    .DE(_00072_),
    .Q(\w[53][16] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][17]$_SDFFCE_PN0P_  (.D(_02226_),
    .DE(_00072_),
    .Q(\w[53][17] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][18]$_SDFFCE_PN0P_  (.D(_02227_),
    .DE(_00072_),
    .Q(\w[53][18] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][19]$_SDFFCE_PN0P_  (.D(_02228_),
    .DE(_00072_),
    .Q(\w[53][19] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][1]$_SDFFCE_PN0P_  (.D(_02229_),
    .DE(_00072_),
    .Q(\w[53][1] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][20]$_SDFFCE_PN0P_  (.D(_02230_),
    .DE(_00072_),
    .Q(\w[53][20] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][21]$_SDFFCE_PN0P_  (.D(_02231_),
    .DE(_00072_),
    .Q(\w[53][21] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][22]$_SDFFCE_PN0P_  (.D(_02232_),
    .DE(_00072_),
    .Q(\w[53][22] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][23]$_SDFFCE_PN0P_  (.D(_02233_),
    .DE(_00072_),
    .Q(\w[53][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][24]$_SDFFCE_PN0P_  (.D(_02234_),
    .DE(_00072_),
    .Q(\w[53][24] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][25]$_SDFFCE_PN0P_  (.D(_02235_),
    .DE(_00072_),
    .Q(\w[53][25] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][26]$_SDFFCE_PN0P_  (.D(_02236_),
    .DE(_00072_),
    .Q(\w[53][26] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][27]$_SDFFCE_PN0P_  (.D(_02237_),
    .DE(_00072_),
    .Q(\w[53][27] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][28]$_SDFFCE_PN0P_  (.D(_02238_),
    .DE(_00072_),
    .Q(\w[53][28] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][29]$_SDFFCE_PN0P_  (.D(_02239_),
    .DE(_00072_),
    .Q(\w[53][29] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][2]$_SDFFCE_PN0P_  (.D(_02240_),
    .DE(_00072_),
    .Q(\w[53][2] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][30]$_SDFFCE_PN0P_  (.D(_02241_),
    .DE(_00072_),
    .Q(\w[53][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][31]$_SDFFCE_PN0P_  (.D(_02242_),
    .DE(_00072_),
    .Q(\w[53][31] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][3]$_SDFFCE_PN0P_  (.D(_02243_),
    .DE(_00072_),
    .Q(\w[53][3] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][4]$_SDFFCE_PN0P_  (.D(_02244_),
    .DE(_00072_),
    .Q(\w[53][4] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][5]$_SDFFCE_PN0P_  (.D(_02245_),
    .DE(_00072_),
    .Q(\w[53][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][6]$_SDFFCE_PN0P_  (.D(_02246_),
    .DE(_00072_),
    .Q(\w[53][6] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][7]$_SDFFCE_PN0P_  (.D(_02247_),
    .DE(_00072_),
    .Q(\w[53][7] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][8]$_SDFFCE_PN0P_  (.D(_02248_),
    .DE(_00072_),
    .Q(\w[53][8] ),
    .CLK(clknet_leaf_252_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[53][9]$_SDFFCE_PN0P_  (.D(_02249_),
    .DE(_00072_),
    .Q(\w[53][9] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][0]$_SDFFCE_PN0P_  (.D(_02250_),
    .DE(_00102_),
    .Q(\w[54][0] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][10]$_SDFFCE_PN0P_  (.D(_02251_),
    .DE(_00102_),
    .Q(\w[54][10] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][11]$_SDFFCE_PN0P_  (.D(_02252_),
    .DE(_00102_),
    .Q(\w[54][11] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][12]$_SDFFCE_PN0P_  (.D(_02253_),
    .DE(_00102_),
    .Q(\w[54][12] ),
    .CLK(clknet_leaf_47_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][13]$_SDFFCE_PN0P_  (.D(_02254_),
    .DE(_00102_),
    .Q(\w[54][13] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][14]$_SDFFCE_PN0P_  (.D(_02255_),
    .DE(_00102_),
    .Q(\w[54][14] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][15]$_SDFFCE_PN0P_  (.D(_02256_),
    .DE(_00102_),
    .Q(\w[54][15] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][16]$_SDFFCE_PN0P_  (.D(_02257_),
    .DE(_00102_),
    .Q(\w[54][16] ),
    .CLK(clknet_leaf_42_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][17]$_SDFFCE_PN0P_  (.D(_02258_),
    .DE(_00102_),
    .Q(\w[54][17] ),
    .CLK(clknet_leaf_110_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][18]$_SDFFCE_PN0P_  (.D(_02259_),
    .DE(_00102_),
    .Q(\w[54][18] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][19]$_SDFFCE_PN0P_  (.D(_02260_),
    .DE(_00102_),
    .Q(\w[54][19] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][1]$_SDFFCE_PN0P_  (.D(_02261_),
    .DE(_00102_),
    .Q(\w[54][1] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][20]$_SDFFCE_PN0P_  (.D(_02262_),
    .DE(_00102_),
    .Q(\w[54][20] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][21]$_SDFFCE_PN0P_  (.D(_02263_),
    .DE(_00102_),
    .Q(\w[54][21] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][22]$_SDFFCE_PN0P_  (.D(_02264_),
    .DE(_00102_),
    .Q(\w[54][22] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][23]$_SDFFCE_PN0P_  (.D(_02265_),
    .DE(_00102_),
    .Q(\w[54][23] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][24]$_SDFFCE_PN0P_  (.D(_02266_),
    .DE(_00102_),
    .Q(\w[54][24] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][25]$_SDFFCE_PN0P_  (.D(_02267_),
    .DE(_00102_),
    .Q(\w[54][25] ),
    .CLK(clknet_leaf_115_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][26]$_SDFFCE_PN0P_  (.D(_02268_),
    .DE(_00102_),
    .Q(\w[54][26] ),
    .CLK(clknet_leaf_108_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][27]$_SDFFCE_PN0P_  (.D(_02269_),
    .DE(_00102_),
    .Q(\w[54][27] ),
    .CLK(clknet_leaf_84_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][28]$_SDFFCE_PN0P_  (.D(_02270_),
    .DE(_00102_),
    .Q(\w[54][28] ),
    .CLK(clknet_leaf_87_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][29]$_SDFFCE_PN0P_  (.D(_02271_),
    .DE(_00102_),
    .Q(\w[54][29] ),
    .CLK(clknet_leaf_70_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][2]$_SDFFCE_PN0P_  (.D(_02272_),
    .DE(_00102_),
    .Q(\w[54][2] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][30]$_SDFFCE_PN0P_  (.D(_02273_),
    .DE(_00102_),
    .Q(\w[54][30] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][31]$_SDFFCE_PN0P_  (.D(_02274_),
    .DE(_00102_),
    .Q(\w[54][31] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][3]$_SDFFCE_PN0P_  (.D(_02275_),
    .DE(_00102_),
    .Q(\w[54][3] ),
    .CLK(clknet_leaf_53_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][4]$_SDFFCE_PN0P_  (.D(_02276_),
    .DE(_00102_),
    .Q(\w[54][4] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][5]$_SDFFCE_PN0P_  (.D(_02277_),
    .DE(_00102_),
    .Q(\w[54][5] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][6]$_SDFFCE_PN0P_  (.D(_02278_),
    .DE(_00102_),
    .Q(\w[54][6] ),
    .CLK(clknet_leaf_50_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][7]$_SDFFCE_PN0P_  (.D(_02279_),
    .DE(_00102_),
    .Q(\w[54][7] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][8]$_SDFFCE_PN0P_  (.D(_02280_),
    .DE(_00102_),
    .Q(\w[54][8] ),
    .CLK(clknet_leaf_106_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[54][9]$_SDFFCE_PN0P_  (.D(_02281_),
    .DE(_00102_),
    .Q(\w[54][9] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][0]$_SDFFCE_PN0P_  (.D(_02282_),
    .DE(net296),
    .Q(\w[55][0] ),
    .CLK(clknet_leaf_278_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][10]$_SDFFCE_PN0P_  (.D(_02283_),
    .DE(net297),
    .Q(\w[55][10] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][11]$_SDFFCE_PN0P_  (.D(_02284_),
    .DE(net297),
    .Q(\w[55][11] ),
    .CLK(clknet_leaf_39_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][12]$_SDFFCE_PN0P_  (.D(_02285_),
    .DE(net297),
    .Q(\w[55][12] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][13]$_SDFFCE_PN0P_  (.D(_02286_),
    .DE(net297),
    .Q(\w[55][13] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][14]$_SDFFCE_PN0P_  (.D(_02287_),
    .DE(net296),
    .Q(\w[55][14] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][15]$_SDFFCE_PN0P_  (.D(_02288_),
    .DE(_00071_),
    .Q(\w[55][15] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][16]$_SDFFCE_PN0P_  (.D(_02289_),
    .DE(net296),
    .Q(\w[55][16] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][17]$_SDFFCE_PN0P_  (.D(_02290_),
    .DE(net296),
    .Q(\w[55][17] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][18]$_SDFFCE_PN0P_  (.D(_02291_),
    .DE(net297),
    .Q(\w[55][18] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][19]$_SDFFCE_PN0P_  (.D(_02292_),
    .DE(net297),
    .Q(\w[55][19] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][1]$_SDFFCE_PN0P_  (.D(_02293_),
    .DE(net296),
    .Q(\w[55][1] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][20]$_SDFFCE_PN0P_  (.D(_02294_),
    .DE(net297),
    .Q(\w[55][20] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][21]$_SDFFCE_PN0P_  (.D(_02295_),
    .DE(net297),
    .Q(\w[55][21] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][22]$_SDFFCE_PN0P_  (.D(_02296_),
    .DE(net297),
    .Q(\w[55][22] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][23]$_SDFFCE_PN0P_  (.D(_02297_),
    .DE(_00071_),
    .Q(\w[55][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][24]$_SDFFCE_PN0P_  (.D(_02298_),
    .DE(net296),
    .Q(\w[55][24] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][25]$_SDFFCE_PN0P_  (.D(_02299_),
    .DE(net296),
    .Q(\w[55][25] ),
    .CLK(clknet_leaf_263_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][26]$_SDFFCE_PN0P_  (.D(_02300_),
    .DE(_00071_),
    .Q(\w[55][26] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][27]$_SDFFCE_PN0P_  (.D(_02301_),
    .DE(net296),
    .Q(\w[55][27] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][28]$_SDFFCE_PN0P_  (.D(_02302_),
    .DE(_00071_),
    .Q(\w[55][28] ),
    .CLK(clknet_leaf_14_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][29]$_SDFFCE_PN0P_  (.D(_02303_),
    .DE(_00071_),
    .Q(\w[55][29] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][2]$_SDFFCE_PN0P_  (.D(_02304_),
    .DE(net296),
    .Q(\w[55][2] ),
    .CLK(clknet_leaf_276_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][30]$_SDFFCE_PN0P_  (.D(_02305_),
    .DE(net297),
    .Q(\w[55][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][31]$_SDFFCE_PN0P_  (.D(_02306_),
    .DE(_00071_),
    .Q(\w[55][31] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][3]$_SDFFCE_PN0P_  (.D(_02307_),
    .DE(_00071_),
    .Q(\w[55][3] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][4]$_SDFFCE_PN0P_  (.D(_02308_),
    .DE(net296),
    .Q(\w[55][4] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][5]$_SDFFCE_PN0P_  (.D(_02309_),
    .DE(_00071_),
    .Q(\w[55][5] ),
    .CLK(clknet_leaf_6_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][6]$_SDFFCE_PN0P_  (.D(_02310_),
    .DE(net296),
    .Q(\w[55][6] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][7]$_SDFFCE_PN0P_  (.D(_02311_),
    .DE(_00071_),
    .Q(\w[55][7] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][8]$_SDFFCE_PN0P_  (.D(_02312_),
    .DE(net296),
    .Q(\w[55][8] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[55][9]$_SDFFCE_PN0P_  (.D(_02313_),
    .DE(_00071_),
    .Q(\w[55][9] ),
    .CLK(clknet_leaf_32_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][0]$_SDFFCE_PN0P_  (.D(_02314_),
    .DE(_00101_),
    .Q(\w[56][0] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][10]$_SDFFCE_PN0P_  (.D(_02315_),
    .DE(_00101_),
    .Q(\w[56][10] ),
    .CLK(clknet_leaf_123_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][11]$_SDFFCE_PN0P_  (.D(_02316_),
    .DE(_00101_),
    .Q(\w[56][11] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][12]$_SDFFCE_PN0P_  (.D(_02317_),
    .DE(_00101_),
    .Q(\w[56][12] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][13]$_SDFFCE_PN0P_  (.D(_02318_),
    .DE(_00101_),
    .Q(\w[56][13] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][14]$_SDFFCE_PN0P_  (.D(_02319_),
    .DE(_00101_),
    .Q(\w[56][14] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][15]$_SDFFCE_PN0P_  (.D(_02320_),
    .DE(_00101_),
    .Q(\w[56][15] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][16]$_SDFFCE_PN0P_  (.D(_02321_),
    .DE(_00101_),
    .Q(\w[56][16] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][17]$_SDFFCE_PN0P_  (.D(_02322_),
    .DE(_00101_),
    .Q(\w[56][17] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][18]$_SDFFCE_PN0P_  (.D(_02323_),
    .DE(_00101_),
    .Q(\w[56][18] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][19]$_SDFFCE_PN0P_  (.D(_02324_),
    .DE(_00101_),
    .Q(\w[56][19] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][1]$_SDFFCE_PN0P_  (.D(_02325_),
    .DE(_00101_),
    .Q(\w[56][1] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][20]$_SDFFCE_PN0P_  (.D(_02326_),
    .DE(_00101_),
    .Q(\w[56][20] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][21]$_SDFFCE_PN0P_  (.D(_02327_),
    .DE(_00101_),
    .Q(\w[56][21] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][22]$_SDFFCE_PN0P_  (.D(_02328_),
    .DE(_00101_),
    .Q(\w[56][22] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][23]$_SDFFCE_PN0P_  (.D(_02329_),
    .DE(_00101_),
    .Q(\w[56][23] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][24]$_SDFFCE_PN0P_  (.D(_02330_),
    .DE(_00101_),
    .Q(\w[56][24] ),
    .CLK(clknet_leaf_140_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][25]$_SDFFCE_PN0P_  (.D(_02331_),
    .DE(_00101_),
    .Q(\w[56][25] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][26]$_SDFFCE_PN0P_  (.D(_02332_),
    .DE(_00101_),
    .Q(\w[56][26] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][27]$_SDFFCE_PN0P_  (.D(_02333_),
    .DE(_00101_),
    .Q(\w[56][27] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][28]$_SDFFCE_PN0P_  (.D(_02334_),
    .DE(_00101_),
    .Q(\w[56][28] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][29]$_SDFFCE_PN0P_  (.D(_02335_),
    .DE(_00101_),
    .Q(\w[56][29] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][2]$_SDFFCE_PN0P_  (.D(_02336_),
    .DE(_00101_),
    .Q(\w[56][2] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][30]$_SDFFCE_PN0P_  (.D(_02337_),
    .DE(_00101_),
    .Q(\w[56][30] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][31]$_SDFFCE_PN0P_  (.D(_02338_),
    .DE(_00101_),
    .Q(\w[56][31] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][3]$_SDFFCE_PN0P_  (.D(_02339_),
    .DE(_00101_),
    .Q(\w[56][3] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][4]$_SDFFCE_PN0P_  (.D(_02340_),
    .DE(_00101_),
    .Q(\w[56][4] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][5]$_SDFFCE_PN0P_  (.D(_02341_),
    .DE(_00101_),
    .Q(\w[56][5] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][6]$_SDFFCE_PN0P_  (.D(_02342_),
    .DE(_00101_),
    .Q(\w[56][6] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][7]$_SDFFCE_PN0P_  (.D(_02343_),
    .DE(_00101_),
    .Q(\w[56][7] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][8]$_SDFFCE_PN0P_  (.D(_02344_),
    .DE(_00101_),
    .Q(\w[56][8] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[56][9]$_SDFFCE_PN0P_  (.D(_02345_),
    .DE(_00101_),
    .Q(\w[56][9] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][0]$_SDFFCE_PN0P_  (.D(_02346_),
    .DE(_00070_),
    .Q(\w[57][0] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][10]$_SDFFCE_PN0P_  (.D(_02347_),
    .DE(_00070_),
    .Q(\w[57][10] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][11]$_SDFFCE_PN0P_  (.D(_02348_),
    .DE(_00070_),
    .Q(\w[57][11] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][12]$_SDFFCE_PN0P_  (.D(_02349_),
    .DE(_00070_),
    .Q(\w[57][12] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][13]$_SDFFCE_PN0P_  (.D(_02350_),
    .DE(_00070_),
    .Q(\w[57][13] ),
    .CLK(clknet_leaf_244_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][14]$_SDFFCE_PN0P_  (.D(_02351_),
    .DE(_00070_),
    .Q(\w[57][14] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][15]$_SDFFCE_PN0P_  (.D(_02352_),
    .DE(_00070_),
    .Q(\w[57][15] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][16]$_SDFFCE_PN0P_  (.D(_02353_),
    .DE(_00070_),
    .Q(\w[57][16] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][17]$_SDFFCE_PN0P_  (.D(_02354_),
    .DE(_00070_),
    .Q(\w[57][17] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][18]$_SDFFCE_PN0P_  (.D(_02355_),
    .DE(_00070_),
    .Q(\w[57][18] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][19]$_SDFFCE_PN0P_  (.D(_02356_),
    .DE(_00070_),
    .Q(\w[57][19] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][1]$_SDFFCE_PN0P_  (.D(_02357_),
    .DE(_00070_),
    .Q(\w[57][1] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][20]$_SDFFCE_PN0P_  (.D(_02358_),
    .DE(_00070_),
    .Q(\w[57][20] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][21]$_SDFFCE_PN0P_  (.D(_02359_),
    .DE(_00070_),
    .Q(\w[57][21] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][22]$_SDFFCE_PN0P_  (.D(_02360_),
    .DE(_00070_),
    .Q(\w[57][22] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][23]$_SDFFCE_PN0P_  (.D(_02361_),
    .DE(_00070_),
    .Q(\w[57][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][24]$_SDFFCE_PN0P_  (.D(_02362_),
    .DE(_00070_),
    .Q(\w[57][24] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][25]$_SDFFCE_PN0P_  (.D(_02363_),
    .DE(_00070_),
    .Q(\w[57][25] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][26]$_SDFFCE_PN0P_  (.D(_02364_),
    .DE(_00070_),
    .Q(\w[57][26] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][27]$_SDFFCE_PN0P_  (.D(_02365_),
    .DE(_00070_),
    .Q(\w[57][27] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][28]$_SDFFCE_PN0P_  (.D(_02366_),
    .DE(_00070_),
    .Q(\w[57][28] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][29]$_SDFFCE_PN0P_  (.D(_02367_),
    .DE(_00070_),
    .Q(\w[57][29] ),
    .CLK(clknet_leaf_28_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][2]$_SDFFCE_PN0P_  (.D(_02368_),
    .DE(_00070_),
    .Q(\w[57][2] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][30]$_SDFFCE_PN0P_  (.D(_02369_),
    .DE(_00070_),
    .Q(\w[57][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][31]$_SDFFCE_PN0P_  (.D(_02370_),
    .DE(_00070_),
    .Q(\w[57][31] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][3]$_SDFFCE_PN0P_  (.D(_02371_),
    .DE(_00070_),
    .Q(\w[57][3] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][4]$_SDFFCE_PN0P_  (.D(_02372_),
    .DE(_00070_),
    .Q(\w[57][4] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][5]$_SDFFCE_PN0P_  (.D(_02373_),
    .DE(_00070_),
    .Q(\w[57][5] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][6]$_SDFFCE_PN0P_  (.D(_02374_),
    .DE(_00070_),
    .Q(\w[57][6] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][7]$_SDFFCE_PN0P_  (.D(_02375_),
    .DE(_00070_),
    .Q(\w[57][7] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][8]$_SDFFCE_PN0P_  (.D(_02376_),
    .DE(_00070_),
    .Q(\w[57][8] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[57][9]$_SDFFCE_PN0P_  (.D(_02377_),
    .DE(_00070_),
    .Q(\w[57][9] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][0]$_SDFFCE_PN0P_  (.D(_02378_),
    .DE(_00100_),
    .Q(\w[58][0] ),
    .CLK(clknet_leaf_128_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][10]$_SDFFCE_PN0P_  (.D(_02379_),
    .DE(_00100_),
    .Q(\w[58][10] ),
    .CLK(clknet_leaf_125_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][11]$_SDFFCE_PN0P_  (.D(_02380_),
    .DE(_00100_),
    .Q(\w[58][11] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][12]$_SDFFCE_PN0P_  (.D(_02381_),
    .DE(_00100_),
    .Q(\w[58][12] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][13]$_SDFFCE_PN0P_  (.D(_02382_),
    .DE(_00100_),
    .Q(\w[58][13] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][14]$_SDFFCE_PN0P_  (.D(_02383_),
    .DE(_00100_),
    .Q(\w[58][14] ),
    .CLK(clknet_leaf_44_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][15]$_SDFFCE_PN0P_  (.D(_02384_),
    .DE(_00100_),
    .Q(\w[58][15] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][16]$_SDFFCE_PN0P_  (.D(_02385_),
    .DE(_00100_),
    .Q(\w[58][16] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][17]$_SDFFCE_PN0P_  (.D(_02386_),
    .DE(_00100_),
    .Q(\w[58][17] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][18]$_SDFFCE_PN0P_  (.D(_02387_),
    .DE(_00100_),
    .Q(\w[58][18] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][19]$_SDFFCE_PN0P_  (.D(_02388_),
    .DE(_00100_),
    .Q(\w[58][19] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][1]$_SDFFCE_PN0P_  (.D(_02389_),
    .DE(_00100_),
    .Q(\w[58][1] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][20]$_SDFFCE_PN0P_  (.D(_02390_),
    .DE(_00100_),
    .Q(\w[58][20] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][21]$_SDFFCE_PN0P_  (.D(_02391_),
    .DE(_00100_),
    .Q(\w[58][21] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][22]$_SDFFCE_PN0P_  (.D(_02392_),
    .DE(_00100_),
    .Q(\w[58][22] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][23]$_SDFFCE_PN0P_  (.D(_02393_),
    .DE(_00100_),
    .Q(\w[58][23] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][24]$_SDFFCE_PN0P_  (.D(_02394_),
    .DE(_00100_),
    .Q(\w[58][24] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][25]$_SDFFCE_PN0P_  (.D(_02395_),
    .DE(_00100_),
    .Q(\w[58][25] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][26]$_SDFFCE_PN0P_  (.D(_02396_),
    .DE(_00100_),
    .Q(\w[58][26] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][27]$_SDFFCE_PN0P_  (.D(_02397_),
    .DE(_00100_),
    .Q(\w[58][27] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][28]$_SDFFCE_PN0P_  (.D(_02398_),
    .DE(_00100_),
    .Q(\w[58][28] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][29]$_SDFFCE_PN0P_  (.D(_02399_),
    .DE(_00100_),
    .Q(\w[58][29] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][2]$_SDFFCE_PN0P_  (.D(_02400_),
    .DE(_00100_),
    .Q(\w[58][2] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][30]$_SDFFCE_PN0P_  (.D(_02401_),
    .DE(_00100_),
    .Q(\w[58][30] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][31]$_SDFFCE_PN0P_  (.D(_02402_),
    .DE(_00100_),
    .Q(\w[58][31] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][3]$_SDFFCE_PN0P_  (.D(_02403_),
    .DE(_00100_),
    .Q(\w[58][3] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][4]$_SDFFCE_PN0P_  (.D(_02404_),
    .DE(_00100_),
    .Q(\w[58][4] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][5]$_SDFFCE_PN0P_  (.D(_02405_),
    .DE(_00100_),
    .Q(\w[58][5] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][6]$_SDFFCE_PN0P_  (.D(_02406_),
    .DE(_00100_),
    .Q(\w[58][6] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][7]$_SDFFCE_PN0P_  (.D(_02407_),
    .DE(_00100_),
    .Q(\w[58][7] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][8]$_SDFFCE_PN0P_  (.D(_02408_),
    .DE(_00100_),
    .Q(\w[58][8] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[58][9]$_SDFFCE_PN0P_  (.D(_02409_),
    .DE(_00100_),
    .Q(\w[58][9] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][0]$_SDFFCE_PN0P_  (.D(_02410_),
    .DE(_00069_),
    .Q(\w[59][0] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][10]$_SDFFCE_PN0P_  (.D(_02411_),
    .DE(_00069_),
    .Q(\w[59][10] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][11]$_SDFFCE_PN0P_  (.D(_02412_),
    .DE(_00069_),
    .Q(\w[59][11] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][12]$_SDFFCE_PN0P_  (.D(_02413_),
    .DE(_00069_),
    .Q(\w[59][12] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][13]$_SDFFCE_PN0P_  (.D(_02414_),
    .DE(_00069_),
    .Q(\w[59][13] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][14]$_SDFFCE_PN0P_  (.D(_02415_),
    .DE(_00069_),
    .Q(\w[59][14] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][15]$_SDFFCE_PN0P_  (.D(_02416_),
    .DE(_00069_),
    .Q(\w[59][15] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][16]$_SDFFCE_PN0P_  (.D(_02417_),
    .DE(_00069_),
    .Q(\w[59][16] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][17]$_SDFFCE_PN0P_  (.D(_02418_),
    .DE(_00069_),
    .Q(\w[59][17] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][18]$_SDFFCE_PN0P_  (.D(_02419_),
    .DE(_00069_),
    .Q(\w[59][18] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][19]$_SDFFCE_PN0P_  (.D(_02420_),
    .DE(_00069_),
    .Q(\w[59][19] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][1]$_SDFFCE_PN0P_  (.D(_02421_),
    .DE(_00069_),
    .Q(\w[59][1] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][20]$_SDFFCE_PN0P_  (.D(_02422_),
    .DE(_00069_),
    .Q(\w[59][20] ),
    .CLK(clknet_leaf_246_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][21]$_SDFFCE_PN0P_  (.D(_02423_),
    .DE(_00069_),
    .Q(\w[59][21] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][22]$_SDFFCE_PN0P_  (.D(_02424_),
    .DE(_00069_),
    .Q(\w[59][22] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][23]$_SDFFCE_PN0P_  (.D(_02425_),
    .DE(_00069_),
    .Q(\w[59][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][24]$_SDFFCE_PN0P_  (.D(_02426_),
    .DE(_00069_),
    .Q(\w[59][24] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][25]$_SDFFCE_PN0P_  (.D(_02427_),
    .DE(_00069_),
    .Q(\w[59][25] ),
    .CLK(clknet_leaf_262_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][26]$_SDFFCE_PN0P_  (.D(_02428_),
    .DE(_00069_),
    .Q(\w[59][26] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][27]$_SDFFCE_PN0P_  (.D(_02429_),
    .DE(_00069_),
    .Q(\w[59][27] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][28]$_SDFFCE_PN0P_  (.D(_02430_),
    .DE(_00069_),
    .Q(\w[59][28] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][29]$_SDFFCE_PN0P_  (.D(_02431_),
    .DE(_00069_),
    .Q(\w[59][29] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][2]$_SDFFCE_PN0P_  (.D(_02432_),
    .DE(_00069_),
    .Q(\w[59][2] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][30]$_SDFFCE_PN0P_  (.D(_02433_),
    .DE(_00069_),
    .Q(\w[59][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][31]$_SDFFCE_PN0P_  (.D(_02434_),
    .DE(_00069_),
    .Q(\w[59][31] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][3]$_SDFFCE_PN0P_  (.D(_02435_),
    .DE(_00069_),
    .Q(\w[59][3] ),
    .CLK(clknet_leaf_4_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][4]$_SDFFCE_PN0P_  (.D(_02436_),
    .DE(_00069_),
    .Q(\w[59][4] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][5]$_SDFFCE_PN0P_  (.D(_02437_),
    .DE(_00069_),
    .Q(\w[59][5] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][6]$_SDFFCE_PN0P_  (.D(_02438_),
    .DE(_00069_),
    .Q(\w[59][6] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][7]$_SDFFCE_PN0P_  (.D(_02439_),
    .DE(_00069_),
    .Q(\w[59][7] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][8]$_SDFFCE_PN0P_  (.D(_02440_),
    .DE(_00069_),
    .Q(\w[59][8] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[59][9]$_SDFFCE_PN0P_  (.D(_02441_),
    .DE(_00069_),
    .Q(\w[59][9] ),
    .CLK(clknet_leaf_36_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][0]$_DFFE_PP_  (.D(_00481_),
    .DE(_00068_),
    .Q(\w[5][0] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][10]$_DFFE_PP_  (.D(_00482_),
    .DE(_00068_),
    .Q(\w[5][10] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][11]$_DFFE_PP_  (.D(_00483_),
    .DE(_00068_),
    .Q(\w[5][11] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][12]$_DFFE_PP_  (.D(_00484_),
    .DE(_00068_),
    .Q(\w[5][12] ),
    .CLK(clknet_leaf_222_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][13]$_DFFE_PP_  (.D(_00485_),
    .DE(_00068_),
    .Q(\w[5][13] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][14]$_DFFE_PP_  (.D(_00486_),
    .DE(_00068_),
    .Q(\w[5][14] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][15]$_DFFE_PP_  (.D(_00487_),
    .DE(_00068_),
    .Q(\w[5][15] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][16]$_DFFE_PP_  (.D(_00488_),
    .DE(_00068_),
    .Q(\w[5][16] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][17]$_DFFE_PP_  (.D(_00489_),
    .DE(_00068_),
    .Q(\w[5][17] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][18]$_DFFE_PP_  (.D(_00490_),
    .DE(_00068_),
    .Q(\w[5][18] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][19]$_DFFE_PP_  (.D(_00491_),
    .DE(_00068_),
    .Q(\w[5][19] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][1]$_DFFE_PP_  (.D(_00492_),
    .DE(_00068_),
    .Q(\w[5][1] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][20]$_DFFE_PP_  (.D(_00493_),
    .DE(_00068_),
    .Q(\w[5][20] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][21]$_DFFE_PP_  (.D(_00494_),
    .DE(_00068_),
    .Q(\w[5][21] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][22]$_DFFE_PP_  (.D(_00495_),
    .DE(_00068_),
    .Q(\w[5][22] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][23]$_DFFE_PP_  (.D(_00496_),
    .DE(_00068_),
    .Q(\w[5][23] ),
    .CLK(clknet_leaf_19_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][24]$_DFFE_PP_  (.D(_00497_),
    .DE(_00068_),
    .Q(\w[5][24] ),
    .CLK(clknet_leaf_277_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][25]$_DFFE_PP_  (.D(_00498_),
    .DE(_00068_),
    .Q(\w[5][25] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][26]$_DFFE_PP_  (.D(_00499_),
    .DE(_00068_),
    .Q(\w[5][26] ),
    .CLK(clknet_leaf_20_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][27]$_DFFE_PP_  (.D(_00500_),
    .DE(_00068_),
    .Q(\w[5][27] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][28]$_DFFE_PP_  (.D(_00501_),
    .DE(_00068_),
    .Q(\w[5][28] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][29]$_DFFE_PP_  (.D(_00502_),
    .DE(_00068_),
    .Q(\w[5][29] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][2]$_DFFE_PP_  (.D(_00503_),
    .DE(_00068_),
    .Q(\w[5][2] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][30]$_DFFE_PP_  (.D(_00504_),
    .DE(_00068_),
    .Q(\w[5][30] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][31]$_DFFE_PP_  (.D(_00505_),
    .DE(_00068_),
    .Q(\w[5][31] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][3]$_DFFE_PP_  (.D(_00506_),
    .DE(_00068_),
    .Q(\w[5][3] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][4]$_DFFE_PP_  (.D(_00507_),
    .DE(_00068_),
    .Q(\w[5][4] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][5]$_DFFE_PP_  (.D(_00508_),
    .DE(_00068_),
    .Q(\w[5][5] ),
    .CLK(clknet_leaf_282_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][6]$_DFFE_PP_  (.D(_00509_),
    .DE(_00068_),
    .Q(\w[5][6] ),
    .CLK(clknet_leaf_267_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][7]$_DFFE_PP_  (.D(_00510_),
    .DE(_00068_),
    .Q(\w[5][7] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][8]$_DFFE_PP_  (.D(_00511_),
    .DE(_00068_),
    .Q(\w[5][8] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[5][9]$_DFFE_PP_  (.D(_00512_),
    .DE(_00068_),
    .Q(\w[5][9] ),
    .CLK(clknet_leaf_26_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][0]$_SDFFCE_PN0P_  (.D(_02442_),
    .DE(_00099_),
    .Q(\w[60][0] ),
    .CLK(clknet_leaf_130_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][10]$_SDFFCE_PN0P_  (.D(_02443_),
    .DE(_00099_),
    .Q(\w[60][10] ),
    .CLK(clknet_leaf_124_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][11]$_SDFFCE_PN0P_  (.D(_02444_),
    .DE(_00099_),
    .Q(\w[60][11] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][12]$_SDFFCE_PN0P_  (.D(_02445_),
    .DE(_00099_),
    .Q(\w[60][12] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][13]$_SDFFCE_PN0P_  (.D(_02446_),
    .DE(_00099_),
    .Q(\w[60][13] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][14]$_SDFFCE_PN0P_  (.D(_02447_),
    .DE(_00099_),
    .Q(\w[60][14] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][15]$_SDFFCE_PN0P_  (.D(_02448_),
    .DE(_00099_),
    .Q(\w[60][15] ),
    .CLK(clknet_leaf_54_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][16]$_SDFFCE_PN0P_  (.D(_02449_),
    .DE(_00099_),
    .Q(\w[60][16] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][17]$_SDFFCE_PN0P_  (.D(_02450_),
    .DE(_00099_),
    .Q(\w[60][17] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][18]$_SDFFCE_PN0P_  (.D(_02451_),
    .DE(_00099_),
    .Q(\w[60][18] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][19]$_SDFFCE_PN0P_  (.D(_02452_),
    .DE(_00099_),
    .Q(\w[60][19] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][1]$_SDFFCE_PN0P_  (.D(_02453_),
    .DE(_00099_),
    .Q(\w[60][1] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][20]$_SDFFCE_PN0P_  (.D(_02454_),
    .DE(_00099_),
    .Q(\w[60][20] ),
    .CLK(clknet_leaf_178_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][21]$_SDFFCE_PN0P_  (.D(_02455_),
    .DE(_00099_),
    .Q(\w[60][21] ),
    .CLK(clknet_leaf_120_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][22]$_SDFFCE_PN0P_  (.D(_02456_),
    .DE(_00099_),
    .Q(\w[60][22] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][23]$_SDFFCE_PN0P_  (.D(_02457_),
    .DE(_00099_),
    .Q(\w[60][23] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][24]$_SDFFCE_PN0P_  (.D(_02458_),
    .DE(_00099_),
    .Q(\w[60][24] ),
    .CLK(clknet_leaf_105_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][25]$_SDFFCE_PN0P_  (.D(_02459_),
    .DE(_00099_),
    .Q(\w[60][25] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][26]$_SDFFCE_PN0P_  (.D(_02460_),
    .DE(_00099_),
    .Q(\w[60][26] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][27]$_SDFFCE_PN0P_  (.D(_02461_),
    .DE(_00099_),
    .Q(\w[60][27] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][28]$_SDFFCE_PN0P_  (.D(_02462_),
    .DE(_00099_),
    .Q(\w[60][28] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][29]$_SDFFCE_PN0P_  (.D(_02463_),
    .DE(_00099_),
    .Q(\w[60][29] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][2]$_SDFFCE_PN0P_  (.D(_02464_),
    .DE(_00099_),
    .Q(\w[60][2] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][30]$_SDFFCE_PN0P_  (.D(_02465_),
    .DE(_00099_),
    .Q(\w[60][30] ),
    .CLK(clknet_leaf_71_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][31]$_SDFFCE_PN0P_  (.D(_02466_),
    .DE(_00099_),
    .Q(\w[60][31] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][3]$_SDFFCE_PN0P_  (.D(_02467_),
    .DE(_00099_),
    .Q(\w[60][3] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][4]$_SDFFCE_PN0P_  (.D(_02468_),
    .DE(_00099_),
    .Q(\w[60][4] ),
    .CLK(clknet_leaf_63_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][5]$_SDFFCE_PN0P_  (.D(_02469_),
    .DE(_00099_),
    .Q(\w[60][5] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][6]$_SDFFCE_PN0P_  (.D(_02470_),
    .DE(_00099_),
    .Q(\w[60][6] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][7]$_SDFFCE_PN0P_  (.D(_02471_),
    .DE(_00099_),
    .Q(\w[60][7] ),
    .CLK(clknet_leaf_48_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][8]$_SDFFCE_PN0P_  (.D(_02472_),
    .DE(_00099_),
    .Q(\w[60][8] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[60][9]$_SDFFCE_PN0P_  (.D(_02473_),
    .DE(_00099_),
    .Q(\w[60][9] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][0]$_SDFFCE_PN0P_  (.D(_02474_),
    .DE(_00067_),
    .Q(\w[61][0] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][10]$_SDFFCE_PN0P_  (.D(_02475_),
    .DE(_00067_),
    .Q(\w[61][10] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][11]$_SDFFCE_PN0P_  (.D(_02476_),
    .DE(_00067_),
    .Q(\w[61][11] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][12]$_SDFFCE_PN0P_  (.D(_02477_),
    .DE(_00067_),
    .Q(\w[61][12] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][13]$_SDFFCE_PN0P_  (.D(_02478_),
    .DE(_00067_),
    .Q(\w[61][13] ),
    .CLK(clknet_leaf_245_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][14]$_SDFFCE_PN0P_  (.D(_02479_),
    .DE(_00067_),
    .Q(\w[61][14] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][15]$_SDFFCE_PN0P_  (.D(_02480_),
    .DE(_00067_),
    .Q(\w[61][15] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][16]$_SDFFCE_PN0P_  (.D(_02481_),
    .DE(_00067_),
    .Q(\w[61][16] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][17]$_SDFFCE_PN0P_  (.D(_02482_),
    .DE(_00067_),
    .Q(\w[61][17] ),
    .CLK(clknet_leaf_280_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][18]$_SDFFCE_PN0P_  (.D(_02483_),
    .DE(_00067_),
    .Q(\w[61][18] ),
    .CLK(clknet_leaf_240_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][19]$_SDFFCE_PN0P_  (.D(_02484_),
    .DE(_00067_),
    .Q(\w[61][19] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][1]$_SDFFCE_PN0P_  (.D(_02485_),
    .DE(_00067_),
    .Q(\w[61][1] ),
    .CLK(clknet_leaf_9_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][20]$_SDFFCE_PN0P_  (.D(_02486_),
    .DE(_00067_),
    .Q(\w[61][20] ),
    .CLK(clknet_leaf_179_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][21]$_SDFFCE_PN0P_  (.D(_02487_),
    .DE(_00067_),
    .Q(\w[61][21] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][22]$_SDFFCE_PN0P_  (.D(_02488_),
    .DE(_00067_),
    .Q(\w[61][22] ),
    .CLK(clknet_leaf_228_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][23]$_SDFFCE_PN0P_  (.D(_02489_),
    .DE(_00067_),
    .Q(\w[61][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][24]$_SDFFCE_PN0P_  (.D(_02490_),
    .DE(_00067_),
    .Q(\w[61][24] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][25]$_SDFFCE_PN0P_  (.D(_02491_),
    .DE(_00067_),
    .Q(\w[61][25] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][26]$_SDFFCE_PN0P_  (.D(_02492_),
    .DE(_00067_),
    .Q(\w[61][26] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][27]$_SDFFCE_PN0P_  (.D(_02493_),
    .DE(_00067_),
    .Q(\w[61][27] ),
    .CLK(clknet_leaf_33_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][28]$_SDFFCE_PN0P_  (.D(_02494_),
    .DE(_00067_),
    .Q(\w[61][28] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][29]$_SDFFCE_PN0P_  (.D(_02495_),
    .DE(_00067_),
    .Q(\w[61][29] ),
    .CLK(clknet_leaf_29_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][2]$_SDFFCE_PN0P_  (.D(_02496_),
    .DE(_00067_),
    .Q(\w[61][2] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][30]$_SDFFCE_PN0P_  (.D(_02497_),
    .DE(_00067_),
    .Q(\w[61][30] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][31]$_SDFFCE_PN0P_  (.D(_02498_),
    .DE(_00067_),
    .Q(\w[61][31] ),
    .CLK(clknet_leaf_7_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][3]$_SDFFCE_PN0P_  (.D(_02499_),
    .DE(_00067_),
    .Q(\w[61][3] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][4]$_SDFFCE_PN0P_  (.D(_02500_),
    .DE(_00067_),
    .Q(\w[61][4] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][5]$_SDFFCE_PN0P_  (.D(_02501_),
    .DE(_00067_),
    .Q(\w[61][5] ),
    .CLK(clknet_leaf_5_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][6]$_SDFFCE_PN0P_  (.D(_02502_),
    .DE(_00067_),
    .Q(\w[61][6] ),
    .CLK(clknet_leaf_256_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][7]$_SDFFCE_PN0P_  (.D(_02503_),
    .DE(_00067_),
    .Q(\w[61][7] ),
    .CLK(clknet_leaf_11_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][8]$_SDFFCE_PN0P_  (.D(_02504_),
    .DE(_00067_),
    .Q(\w[61][8] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[61][9]$_SDFFCE_PN0P_  (.D(_02505_),
    .DE(_00067_),
    .Q(\w[61][9] ),
    .CLK(clknet_leaf_35_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][0]$_SDFFCE_PN0P_  (.D(_02506_),
    .DE(_00098_),
    .Q(\w[62][0] ),
    .CLK(clknet_leaf_127_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][10]$_SDFFCE_PN0P_  (.D(_02507_),
    .DE(_00098_),
    .Q(\w[62][10] ),
    .CLK(clknet_leaf_126_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][11]$_SDFFCE_PN0P_  (.D(_02508_),
    .DE(_00098_),
    .Q(\w[62][11] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][12]$_SDFFCE_PN0P_  (.D(_02509_),
    .DE(_00098_),
    .Q(\w[62][12] ),
    .CLK(clknet_leaf_45_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][13]$_SDFFCE_PN0P_  (.D(_02510_),
    .DE(_00098_),
    .Q(\w[62][13] ),
    .CLK(clknet_leaf_43_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][14]$_SDFFCE_PN0P_  (.D(_02511_),
    .DE(_00098_),
    .Q(\w[62][14] ),
    .CLK(clknet_leaf_113_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][15]$_SDFFCE_PN0P_  (.D(_02512_),
    .DE(_00098_),
    .Q(\w[62][15] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][16]$_SDFFCE_PN0P_  (.D(_02513_),
    .DE(_00098_),
    .Q(\w[62][16] ),
    .CLK(clknet_leaf_41_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][17]$_SDFFCE_PN0P_  (.D(_02514_),
    .DE(_00098_),
    .Q(\w[62][17] ),
    .CLK(clknet_leaf_112_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][18]$_SDFFCE_PN0P_  (.D(_02515_),
    .DE(_00098_),
    .Q(\w[62][18] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][19]$_SDFFCE_PN0P_  (.D(_02516_),
    .DE(_00098_),
    .Q(\w[62][19] ),
    .CLK(clknet_leaf_117_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][1]$_SDFFCE_PN0P_  (.D(_02517_),
    .DE(_00098_),
    .Q(\w[62][1] ),
    .CLK(clknet_leaf_122_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][20]$_SDFFCE_PN0P_  (.D(_02518_),
    .DE(_00098_),
    .Q(\w[62][20] ),
    .CLK(clknet_leaf_121_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][21]$_SDFFCE_PN0P_  (.D(_02519_),
    .DE(_00098_),
    .Q(\w[62][21] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][22]$_SDFFCE_PN0P_  (.D(_02520_),
    .DE(_00098_),
    .Q(\w[62][22] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][23]$_SDFFCE_PN0P_  (.D(_02521_),
    .DE(_00098_),
    .Q(\w[62][23] ),
    .CLK(clknet_leaf_111_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][24]$_SDFFCE_PN0P_  (.D(_02522_),
    .DE(_00098_),
    .Q(\w[62][24] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][25]$_SDFFCE_PN0P_  (.D(_02523_),
    .DE(_00098_),
    .Q(\w[62][25] ),
    .CLK(clknet_leaf_114_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][26]$_SDFFCE_PN0P_  (.D(_02524_),
    .DE(_00098_),
    .Q(\w[62][26] ),
    .CLK(clknet_leaf_107_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][27]$_SDFFCE_PN0P_  (.D(_02525_),
    .DE(_00098_),
    .Q(\w[62][27] ),
    .CLK(clknet_leaf_68_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][28]$_SDFFCE_PN0P_  (.D(_02526_),
    .DE(_00098_),
    .Q(\w[62][28] ),
    .CLK(clknet_leaf_86_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][29]$_SDFFCE_PN0P_  (.D(_02527_),
    .DE(_00098_),
    .Q(\w[62][29] ),
    .CLK(clknet_leaf_69_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][2]$_SDFFCE_PN0P_  (.D(_02528_),
    .DE(_00098_),
    .Q(\w[62][2] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][30]$_SDFFCE_PN0P_  (.D(_02529_),
    .DE(_00098_),
    .Q(\w[62][30] ),
    .CLK(clknet_leaf_67_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][31]$_SDFFCE_PN0P_  (.D(_02530_),
    .DE(_00098_),
    .Q(\w[62][31] ),
    .CLK(clknet_leaf_119_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][3]$_SDFFCE_PN0P_  (.D(_02531_),
    .DE(_00098_),
    .Q(\w[62][3] ),
    .CLK(clknet_leaf_52_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][4]$_SDFFCE_PN0P_  (.D(_02532_),
    .DE(_00098_),
    .Q(\w[62][4] ),
    .CLK(clknet_leaf_66_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][5]$_SDFFCE_PN0P_  (.D(_02533_),
    .DE(_00098_),
    .Q(\w[62][5] ),
    .CLK(clknet_leaf_65_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][6]$_SDFFCE_PN0P_  (.D(_02534_),
    .DE(_00098_),
    .Q(\w[62][6] ),
    .CLK(clknet_leaf_51_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][7]$_SDFFCE_PN0P_  (.D(_02535_),
    .DE(_00098_),
    .Q(\w[62][7] ),
    .CLK(clknet_leaf_49_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][8]$_SDFFCE_PN0P_  (.D(_02536_),
    .DE(_00098_),
    .Q(\w[62][8] ),
    .CLK(clknet_leaf_116_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[62][9]$_SDFFCE_PN0P_  (.D(_02537_),
    .DE(_00098_),
    .Q(\w[62][9] ),
    .CLK(clknet_leaf_118_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][0]$_SDFFCE_PN0P_  (.D(_02538_),
    .DE(_00066_),
    .Q(\w[63][0] ),
    .CLK(clknet_leaf_255_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][10]$_SDFFCE_PN0P_  (.D(_02539_),
    .DE(_00066_),
    .Q(\w[63][10] ),
    .CLK(clknet_leaf_250_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][11]$_SDFFCE_PN0P_  (.D(_02540_),
    .DE(_00066_),
    .Q(\w[63][11] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][12]$_SDFFCE_PN0P_  (.D(_02541_),
    .DE(_00066_),
    .Q(\w[63][12] ),
    .CLK(clknet_leaf_248_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][13]$_SDFFCE_PN0P_  (.D(_02542_),
    .DE(_00066_),
    .Q(\w[63][13] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][14]$_SDFFCE_PN0P_  (.D(_02543_),
    .DE(_00066_),
    .Q(\w[63][14] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][15]$_SDFFCE_PN0P_  (.D(_02544_),
    .DE(_00066_),
    .Q(\w[63][15] ),
    .CLK(clknet_leaf_27_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][16]$_SDFFCE_PN0P_  (.D(_02545_),
    .DE(_00066_),
    .Q(\w[63][16] ),
    .CLK(clknet_leaf_253_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][17]$_SDFFCE_PN0P_  (.D(_02546_),
    .DE(_00066_),
    .Q(\w[63][17] ),
    .CLK(clknet_leaf_279_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][18]$_SDFFCE_PN0P_  (.D(_02547_),
    .DE(_00066_),
    .Q(\w[63][18] ),
    .CLK(clknet_leaf_251_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][19]$_SDFFCE_PN0P_  (.D(_02548_),
    .DE(_00066_),
    .Q(\w[63][19] ),
    .CLK(clknet_leaf_247_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][1]$_SDFFCE_PN0P_  (.D(_02549_),
    .DE(_00066_),
    .Q(\w[63][1] ),
    .CLK(clknet_leaf_10_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][20]$_SDFFCE_PN0P_  (.D(_02550_),
    .DE(_00066_),
    .Q(\w[63][20] ),
    .CLK(clknet_leaf_40_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][21]$_SDFFCE_PN0P_  (.D(_02551_),
    .DE(_00066_),
    .Q(\w[63][21] ),
    .CLK(clknet_leaf_260_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][22]$_SDFFCE_PN0P_  (.D(_02552_),
    .DE(_00066_),
    .Q(\w[63][22] ),
    .CLK(clknet_leaf_261_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][23]$_SDFFCE_PN0P_  (.D(_02553_),
    .DE(_00066_),
    .Q(\w[63][23] ),
    .CLK(clknet_leaf_31_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][24]$_SDFFCE_PN0P_  (.D(_02554_),
    .DE(_00066_),
    .Q(\w[63][24] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][25]$_SDFFCE_PN0P_  (.D(_02555_),
    .DE(_00066_),
    .Q(\w[63][25] ),
    .CLK(clknet_leaf_258_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][26]$_SDFFCE_PN0P_  (.D(_02556_),
    .DE(_00066_),
    .Q(\w[63][26] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][27]$_SDFFCE_PN0P_  (.D(_02557_),
    .DE(_00066_),
    .Q(\w[63][27] ),
    .CLK(clknet_leaf_34_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][28]$_SDFFCE_PN0P_  (.D(_02558_),
    .DE(_00066_),
    .Q(\w[63][28] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][29]$_SDFFCE_PN0P_  (.D(_02559_),
    .DE(_00066_),
    .Q(\w[63][29] ),
    .CLK(clknet_leaf_30_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][2]$_SDFFCE_PN0P_  (.D(_02560_),
    .DE(_00066_),
    .Q(\w[63][2] ),
    .CLK(clknet_leaf_257_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][30]$_SDFFCE_PN0P_  (.D(_02561_),
    .DE(_00066_),
    .Q(\w[63][30] ),
    .CLK(clknet_leaf_38_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][31]$_SDFFCE_PN0P_  (.D(_02562_),
    .DE(_00066_),
    .Q(\w[63][31] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][3]$_SDFFCE_PN0P_  (.D(_02563_),
    .DE(_00066_),
    .Q(\w[63][3] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][4]$_SDFFCE_PN0P_  (.D(_02564_),
    .DE(_00066_),
    .Q(\w[63][4] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][5]$_SDFFCE_PN0P_  (.D(_02565_),
    .DE(_00066_),
    .Q(\w[63][5] ),
    .CLK(clknet_leaf_8_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][6]$_SDFFCE_PN0P_  (.D(_02566_),
    .DE(_00066_),
    .Q(\w[63][6] ),
    .CLK(clknet_leaf_254_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][7]$_SDFFCE_PN0P_  (.D(_02567_),
    .DE(_00066_),
    .Q(\w[63][7] ),
    .CLK(clknet_leaf_12_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][8]$_SDFFCE_PN0P_  (.D(_02568_),
    .DE(_00066_),
    .Q(\w[63][8] ),
    .CLK(clknet_leaf_259_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[63][9]$_SDFFCE_PN0P_  (.D(_02569_),
    .DE(_00066_),
    .Q(\w[63][9] ),
    .CLK(clknet_leaf_37_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][0]$_DFFE_PP_  (.D(_00513_),
    .DE(_00097_),
    .Q(\w[6][0] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][10]$_DFFE_PP_  (.D(_00514_),
    .DE(_00097_),
    .Q(\w[6][10] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][11]$_DFFE_PP_  (.D(_00515_),
    .DE(_00097_),
    .Q(\w[6][11] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][12]$_DFFE_PP_  (.D(_00516_),
    .DE(_00097_),
    .Q(\w[6][12] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][13]$_DFFE_PP_  (.D(_00517_),
    .DE(_00097_),
    .Q(\w[6][13] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][14]$_DFFE_PP_  (.D(_00518_),
    .DE(_00097_),
    .Q(\w[6][14] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][15]$_DFFE_PP_  (.D(_00519_),
    .DE(_00097_),
    .Q(\w[6][15] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][16]$_DFFE_PP_  (.D(_00520_),
    .DE(_00097_),
    .Q(\w[6][16] ),
    .CLK(clknet_leaf_59_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][17]$_DFFE_PP_  (.D(_00521_),
    .DE(_00097_),
    .Q(\w[6][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][18]$_DFFE_PP_  (.D(_00522_),
    .DE(_00097_),
    .Q(\w[6][18] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][19]$_DFFE_PP_  (.D(_00523_),
    .DE(_00097_),
    .Q(\w[6][19] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][1]$_DFFE_PP_  (.D(_00524_),
    .DE(_00097_),
    .Q(\w[6][1] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][20]$_DFFE_PP_  (.D(_00525_),
    .DE(_00097_),
    .Q(\w[6][20] ),
    .CLK(clknet_leaf_175_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][21]$_DFFE_PP_  (.D(_00526_),
    .DE(_00097_),
    .Q(\w[6][21] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][22]$_DFFE_PP_  (.D(_00527_),
    .DE(_00097_),
    .Q(\w[6][22] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][23]$_DFFE_PP_  (.D(_00528_),
    .DE(_00097_),
    .Q(\w[6][23] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][24]$_DFFE_PP_  (.D(_00529_),
    .DE(_00097_),
    .Q(\w[6][24] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][25]$_DFFE_PP_  (.D(_00530_),
    .DE(_00097_),
    .Q(\w[6][25] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][26]$_DFFE_PP_  (.D(_00531_),
    .DE(_00097_),
    .Q(\w[6][26] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][27]$_DFFE_PP_  (.D(_00532_),
    .DE(_00097_),
    .Q(\w[6][27] ),
    .CLK(clknet_leaf_81_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][28]$_DFFE_PP_  (.D(_00533_),
    .DE(_00097_),
    .Q(\w[6][28] ),
    .CLK(clknet_leaf_91_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][29]$_DFFE_PP_  (.D(_00534_),
    .DE(_00097_),
    .Q(\w[6][29] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][2]$_DFFE_PP_  (.D(_00535_),
    .DE(_00097_),
    .Q(\w[6][2] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][30]$_DFFE_PP_  (.D(_00536_),
    .DE(_00097_),
    .Q(\w[6][30] ),
    .CLK(clknet_leaf_76_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][31]$_DFFE_PP_  (.D(_00537_),
    .DE(_00097_),
    .Q(\w[6][31] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][3]$_DFFE_PP_  (.D(_00538_),
    .DE(_00097_),
    .Q(\w[6][3] ),
    .CLK(clknet_leaf_58_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][4]$_DFFE_PP_  (.D(_00539_),
    .DE(_00097_),
    .Q(\w[6][4] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][5]$_DFFE_PP_  (.D(_00540_),
    .DE(_00097_),
    .Q(\w[6][5] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][6]$_DFFE_PP_  (.D(_00541_),
    .DE(_00097_),
    .Q(\w[6][6] ),
    .CLK(clknet_leaf_64_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][7]$_DFFE_PP_  (.D(_00542_),
    .DE(_00097_),
    .Q(\w[6][7] ),
    .CLK(clknet_leaf_83_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][8]$_DFFE_PP_  (.D(_00543_),
    .DE(_00097_),
    .Q(\w[6][8] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[6][9]$_DFFE_PP_  (.D(_00544_),
    .DE(_00097_),
    .Q(\w[6][9] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][0]$_DFFE_PP_  (.D(_00545_),
    .DE(_00065_),
    .Q(\w[7][0] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][10]$_DFFE_PP_  (.D(_00546_),
    .DE(_00065_),
    .Q(\w[7][10] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][11]$_DFFE_PP_  (.D(_00547_),
    .DE(_00065_),
    .Q(\w[7][11] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][12]$_DFFE_PP_  (.D(_00548_),
    .DE(_00065_),
    .Q(\w[7][12] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][13]$_DFFE_PP_  (.D(_00549_),
    .DE(_00065_),
    .Q(\w[7][13] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][14]$_DFFE_PP_  (.D(_00550_),
    .DE(_00065_),
    .Q(\w[7][14] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][15]$_DFFE_PP_  (.D(_00551_),
    .DE(_00065_),
    .Q(\w[7][15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][16]$_DFFE_PP_  (.D(_00552_),
    .DE(_00065_),
    .Q(\w[7][16] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][17]$_DFFE_PP_  (.D(_00553_),
    .DE(_00065_),
    .Q(\w[7][17] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][18]$_DFFE_PP_  (.D(_00554_),
    .DE(_00065_),
    .Q(\w[7][18] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][19]$_DFFE_PP_  (.D(_00555_),
    .DE(_00065_),
    .Q(\w[7][19] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][1]$_DFFE_PP_  (.D(_00556_),
    .DE(_00065_),
    .Q(\w[7][1] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][20]$_DFFE_PP_  (.D(_00557_),
    .DE(_00065_),
    .Q(\w[7][20] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][21]$_DFFE_PP_  (.D(_00558_),
    .DE(_00065_),
    .Q(\w[7][21] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][22]$_DFFE_PP_  (.D(_00559_),
    .DE(_00065_),
    .Q(\w[7][22] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][23]$_DFFE_PP_  (.D(_00560_),
    .DE(_00065_),
    .Q(\w[7][23] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][24]$_DFFE_PP_  (.D(_00561_),
    .DE(_00065_),
    .Q(\w[7][24] ),
    .CLK(clknet_leaf_273_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][25]$_DFFE_PP_  (.D(_00562_),
    .DE(_00065_),
    .Q(\w[7][25] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][26]$_DFFE_PP_  (.D(_00563_),
    .DE(_00065_),
    .Q(\w[7][26] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][27]$_DFFE_PP_  (.D(_00564_),
    .DE(_00065_),
    .Q(\w[7][27] ),
    .CLK(clknet_leaf_283_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][28]$_DFFE_PP_  (.D(_00565_),
    .DE(_00065_),
    .Q(\w[7][28] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][29]$_DFFE_PP_  (.D(_00566_),
    .DE(_00065_),
    .Q(\w[7][29] ),
    .CLK(clknet_leaf_22_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][2]$_DFFE_PP_  (.D(_00567_),
    .DE(_00065_),
    .Q(\w[7][2] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][30]$_DFFE_PP_  (.D(_00568_),
    .DE(_00065_),
    .Q(\w[7][30] ),
    .CLK(clknet_leaf_25_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][31]$_DFFE_PP_  (.D(_00569_),
    .DE(_00065_),
    .Q(\w[7][31] ),
    .CLK(clknet_leaf_288_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][3]$_DFFE_PP_  (.D(_00570_),
    .DE(_00065_),
    .Q(\w[7][3] ),
    .CLK(clknet_leaf_281_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][4]$_DFFE_PP_  (.D(_00571_),
    .DE(_00065_),
    .Q(\w[7][4] ),
    .CLK(clknet_leaf_271_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][5]$_DFFE_PP_  (.D(_00572_),
    .DE(_00065_),
    .Q(\w[7][5] ),
    .CLK(clknet_leaf_287_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][6]$_DFFE_PP_  (.D(_00573_),
    .DE(_00065_),
    .Q(\w[7][6] ),
    .CLK(clknet_leaf_269_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][7]$_DFFE_PP_  (.D(_00574_),
    .DE(_00065_),
    .Q(\w[7][7] ),
    .CLK(clknet_leaf_2_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][8]$_DFFE_PP_  (.D(_00575_),
    .DE(_00065_),
    .Q(\w[7][8] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[7][9]$_DFFE_PP_  (.D(_00576_),
    .DE(_00065_),
    .Q(\w[7][9] ),
    .CLK(clknet_leaf_18_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][0]$_DFFE_PP_  (.D(_00577_),
    .DE(_00096_),
    .Q(\w[8][0] ),
    .CLK(clknet_leaf_149_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][10]$_DFFE_PP_  (.D(_00578_),
    .DE(_00096_),
    .Q(\w[8][10] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][11]$_DFFE_PP_  (.D(_00579_),
    .DE(_00096_),
    .Q(\w[8][11] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][12]$_DFFE_PP_  (.D(_00580_),
    .DE(_00096_),
    .Q(\w[8][12] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][13]$_DFFE_PP_  (.D(_00581_),
    .DE(_00096_),
    .Q(\w[8][13] ),
    .CLK(clknet_leaf_89_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][14]$_DFFE_PP_  (.D(_00582_),
    .DE(_00096_),
    .Q(\w[8][14] ),
    .CLK(clknet_leaf_93_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][15]$_DFFE_PP_  (.D(_00583_),
    .DE(_00096_),
    .Q(\w[8][15] ),
    .CLK(clknet_leaf_62_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][16]$_DFFE_PP_  (.D(_00584_),
    .DE(_00096_),
    .Q(\w[8][16] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][17]$_DFFE_PP_  (.D(_00585_),
    .DE(_00096_),
    .Q(\w[8][17] ),
    .CLK(clknet_leaf_94_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][18]$_DFFE_PP_  (.D(_00586_),
    .DE(_00096_),
    .Q(\w[8][18] ),
    .CLK(clknet_leaf_176_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][19]$_DFFE_PP_  (.D(_00587_),
    .DE(_00096_),
    .Q(\w[8][19] ),
    .CLK(clknet_leaf_146_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][1]$_DFFE_PP_  (.D(_00588_),
    .DE(_00096_),
    .Q(\w[8][1] ),
    .CLK(clknet_leaf_145_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][20]$_DFFE_PP_  (.D(_00589_),
    .DE(_00096_),
    .Q(\w[8][20] ),
    .CLK(clknet_leaf_131_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][21]$_DFFE_PP_  (.D(_00590_),
    .DE(_00096_),
    .Q(\w[8][21] ),
    .CLK(clknet_leaf_99_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][22]$_DFFE_PP_  (.D(_00591_),
    .DE(_00096_),
    .Q(\w[8][22] ),
    .CLK(clknet_leaf_147_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][23]$_DFFE_PP_  (.D(_00592_),
    .DE(_00096_),
    .Q(\w[8][23] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][24]$_DFFE_PP_  (.D(_00593_),
    .DE(_00096_),
    .Q(\w[8][24] ),
    .CLK(clknet_leaf_148_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][25]$_DFFE_PP_  (.D(_00594_),
    .DE(_00096_),
    .Q(\w[8][25] ),
    .CLK(clknet_leaf_102_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][26]$_DFFE_PP_  (.D(_00595_),
    .DE(_00096_),
    .Q(\w[8][26] ),
    .CLK(clknet_leaf_98_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][27]$_DFFE_PP_  (.D(_00596_),
    .DE(_00096_),
    .Q(\w[8][27] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][28]$_DFFE_PP_  (.D(_00597_),
    .DE(_00096_),
    .Q(\w[8][28] ),
    .CLK(clknet_leaf_92_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][29]$_DFFE_PP_  (.D(_00598_),
    .DE(_00096_),
    .Q(\w[8][29] ),
    .CLK(clknet_leaf_79_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][2]$_DFFE_PP_  (.D(_00599_),
    .DE(_00096_),
    .Q(\w[8][2] ),
    .CLK(clknet_leaf_80_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][30]$_DFFE_PP_  (.D(_00600_),
    .DE(_00096_),
    .Q(\w[8][30] ),
    .CLK(clknet_leaf_77_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][31]$_DFFE_PP_  (.D(_00601_),
    .DE(_00096_),
    .Q(\w[8][31] ),
    .CLK(clknet_leaf_97_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][3]$_DFFE_PP_  (.D(_00602_),
    .DE(_00096_),
    .Q(\w[8][3] ),
    .CLK(clknet_leaf_57_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][4]$_DFFE_PP_  (.D(_00603_),
    .DE(_00096_),
    .Q(\w[8][4] ),
    .CLK(clknet_leaf_74_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][5]$_DFFE_PP_  (.D(_00604_),
    .DE(_00096_),
    .Q(\w[8][5] ),
    .CLK(clknet_leaf_72_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][6]$_DFFE_PP_  (.D(_00605_),
    .DE(_00096_),
    .Q(\w[8][6] ),
    .CLK(clknet_leaf_60_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][7]$_DFFE_PP_  (.D(_00606_),
    .DE(_00096_),
    .Q(\w[8][7] ),
    .CLK(clknet_leaf_82_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][8]$_DFFE_PP_  (.D(_00607_),
    .DE(_00096_),
    .Q(\w[8][8] ),
    .CLK(clknet_leaf_100_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[8][9]$_DFFE_PP_  (.D(_00608_),
    .DE(_00096_),
    .Q(\w[8][9] ),
    .CLK(clknet_leaf_136_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][0]$_DFFE_PP_  (.D(_00609_),
    .DE(_00064_),
    .Q(\w[9][0] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][10]$_DFFE_PP_  (.D(_00610_),
    .DE(_00064_),
    .Q(\w[9][10] ),
    .CLK(clknet_leaf_237_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][11]$_DFFE_PP_  (.D(_00611_),
    .DE(_00064_),
    .Q(\w[9][11] ),
    .CLK(clknet_leaf_223_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][12]$_DFFE_PP_  (.D(_00612_),
    .DE(_00064_),
    .Q(\w[9][12] ),
    .CLK(clknet_leaf_224_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][13]$_DFFE_PP_  (.D(_00613_),
    .DE(_00064_),
    .Q(\w[9][13] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][14]$_DFFE_PP_  (.D(_00614_),
    .DE(_00064_),
    .Q(\w[9][14] ),
    .CLK(clknet_leaf_268_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][15]$_DFFE_PP_  (.D(_00615_),
    .DE(_00064_),
    .Q(\w[9][15] ),
    .CLK(clknet_leaf_23_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][16]$_DFFE_PP_  (.D(_00616_),
    .DE(_00064_),
    .Q(\w[9][16] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][17]$_DFFE_PP_  (.D(_00617_),
    .DE(_00064_),
    .Q(\w[9][17] ),
    .CLK(clknet_leaf_285_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][18]$_DFFE_PP_  (.D(_00618_),
    .DE(_00064_),
    .Q(\w[9][18] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][19]$_DFFE_PP_  (.D(_00619_),
    .DE(_00064_),
    .Q(\w[9][19] ),
    .CLK(clknet_leaf_238_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][1]$_DFFE_PP_  (.D(_00620_),
    .DE(_00064_),
    .Q(\w[9][1] ),
    .CLK(clknet_leaf_286_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][20]$_DFFE_PP_  (.D(_00621_),
    .DE(_00064_),
    .Q(\w[9][20] ),
    .CLK(clknet_leaf_243_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][21]$_DFFE_PP_  (.D(_00622_),
    .DE(_00064_),
    .Q(\w[9][21] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][22]$_DFFE_PP_  (.D(_00623_),
    .DE(_00064_),
    .Q(\w[9][22] ),
    .CLK(clknet_leaf_221_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][23]$_DFFE_PP_  (.D(_00624_),
    .DE(_00064_),
    .Q(\w[9][23] ),
    .CLK(clknet_leaf_17_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][24]$_DFFE_PP_  (.D(_00625_),
    .DE(_00064_),
    .Q(\w[9][24] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][25]$_DFFE_PP_  (.D(_00626_),
    .DE(_00064_),
    .Q(\w[9][25] ),
    .CLK(clknet_leaf_227_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][26]$_DFFE_PP_  (.D(_00627_),
    .DE(_00064_),
    .Q(\w[9][26] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][27]$_DFFE_PP_  (.D(_00628_),
    .DE(_00064_),
    .Q(\w[9][27] ),
    .CLK(clknet_leaf_284_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][28]$_DFFE_PP_  (.D(_00629_),
    .DE(_00064_),
    .Q(\w[9][28] ),
    .CLK(clknet_leaf_16_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][29]$_DFFE_PP_  (.D(_00630_),
    .DE(_00064_),
    .Q(\w[9][29] ),
    .CLK(clknet_leaf_21_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][2]$_DFFE_PP_  (.D(_00631_),
    .DE(_00064_),
    .Q(\w[9][2] ),
    .CLK(clknet_leaf_270_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][30]$_DFFE_PP_  (.D(_00632_),
    .DE(_00064_),
    .Q(\w[9][30] ),
    .CLK(clknet_leaf_24_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][31]$_DFFE_PP_  (.D(_00633_),
    .DE(_00064_),
    .Q(\w[9][31] ),
    .CLK(clknet_leaf_289_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][3]$_DFFE_PP_  (.D(_00634_),
    .DE(_00064_),
    .Q(\w[9][3] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][4]$_DFFE_PP_  (.D(_00635_),
    .DE(_00064_),
    .Q(\w[9][4] ),
    .CLK(clknet_leaf_272_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][5]$_DFFE_PP_  (.D(_00636_),
    .DE(_00064_),
    .Q(\w[9][5] ),
    .CLK(clknet_leaf_0_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][6]$_DFFE_PP_  (.D(_00637_),
    .DE(_00064_),
    .Q(\w[9][6] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][7]$_DFFE_PP_  (.D(_00638_),
    .DE(_00064_),
    .Q(\w[9][7] ),
    .CLK(clknet_leaf_3_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][8]$_DFFE_PP_  (.D(_00639_),
    .DE(_00064_),
    .Q(\w[9][8] ),
    .CLK(clknet_leaf_266_clk));
 sky130_fd_sc_hd__edfxtp_1 \w[9][9]$_DFFE_PP_  (.D(_00640_),
    .DE(_00064_),
    .Q(\w[9][9] ),
    .CLK(clknet_leaf_13_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[0]$_DFF_P_  (.D(_00000_),
    .Q(\hash.CA1.w_i1[0] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[10]$_DFF_P_  (.D(_00001_),
    .Q(\hash.CA1.w_i1[10] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[11]$_DFF_P_  (.D(_00002_),
    .Q(\hash.CA1.w_i1[11] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[12]$_DFF_P_  (.D(_00003_),
    .Q(\hash.CA1.w_i1[12] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[13]$_DFF_P_  (.D(_00004_),
    .Q(\hash.CA1.w_i1[13] ),
    .CLK(clknet_leaf_139_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[14]$_DFF_P_  (.D(_00005_),
    .Q(\hash.CA1.w_i1[14] ),
    .CLK(clknet_leaf_103_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[15]$_DFF_P_  (.D(_00006_),
    .Q(\hash.CA1.w_i1[15] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[16]$_DFF_P_  (.D(_00007_),
    .Q(\hash.CA1.w_i1[16] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[17]$_DFF_P_  (.D(_00008_),
    .Q(\hash.CA1.w_i1[17] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[18]$_DFF_P_  (.D(_00009_),
    .Q(\hash.CA1.w_i1[18] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[19]$_DFF_P_  (.D(_00010_),
    .Q(\hash.CA1.w_i1[19] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[1]$_DFF_P_  (.D(_00011_),
    .Q(\hash.CA1.w_i1[1] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[20]$_DFF_P_  (.D(_00012_),
    .Q(\hash.CA1.w_i1[20] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[21]$_DFF_P_  (.D(_00013_),
    .Q(\hash.CA1.w_i1[21] ),
    .CLK(clknet_leaf_150_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[22]$_DFF_P_  (.D(_00014_),
    .Q(\hash.CA1.w_i1[22] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[23]$_DFF_P_  (.D(_00015_),
    .Q(\hash.CA1.w_i1[23] ),
    .CLK(clknet_leaf_109_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[24]$_DFF_P_  (.D(_00016_),
    .Q(\hash.CA1.w_i1[24] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[25]$_DFF_P_  (.D(_00017_),
    .Q(\hash.CA1.w_i1[25] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[26]$_DFF_P_  (.D(_00018_),
    .Q(\hash.CA1.w_i1[26] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[27]$_DFF_P_  (.D(_00019_),
    .Q(\hash.CA1.w_i1[27] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[28]$_DFF_P_  (.D(_00020_),
    .Q(\hash.CA1.w_i1[28] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[29]$_DFF_P_  (.D(_00021_),
    .Q(\hash.CA1.w_i1[29] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[2]$_DFF_P_  (.D(_00022_),
    .Q(\hash.CA1.w_i1[2] ),
    .CLK(clknet_leaf_104_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[30]$_DFF_P_  (.D(_00023_),
    .Q(\hash.CA1.w_i1[30] ),
    .CLK(clknet_leaf_152_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[31]$_DFF_P_  (.D(_00024_),
    .Q(\hash.CA1.w_i1[31] ),
    .CLK(clknet_leaf_153_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[3]$_DFF_P_  (.D(_00025_),
    .Q(\hash.CA1.w_i1[3] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[4]$_DFF_P_  (.D(_00026_),
    .Q(\hash.CA1.w_i1[4] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[5]$_DFF_P_  (.D(_00027_),
    .Q(\hash.CA1.w_i1[5] ),
    .CLK(clknet_leaf_133_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[6]$_DFF_P_  (.D(_00028_),
    .Q(\hash.CA1.w_i1[6] ),
    .CLK(clknet_leaf_132_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[7]$_DFF_P_  (.D(_00029_),
    .Q(\hash.CA1.w_i1[7] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[8]$_DFF_P_  (.D(_00030_),
    .Q(\hash.CA1.w_i1[8] ),
    .CLK(clknet_leaf_141_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value1[9]$_DFF_P_  (.D(_00031_),
    .Q(\hash.CA1.w_i1[9] ),
    .CLK(clknet_leaf_135_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[0]$_DFF_P_  (.D(_00032_),
    .Q(\hash.CA1.w_i2[0] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[10]$_DFF_P_  (.D(_00033_),
    .Q(\hash.CA1.w_i2[10] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[11]$_DFF_P_  (.D(_00034_),
    .Q(\hash.CA1.w_i2[11] ),
    .CLK(clknet_leaf_239_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[12]$_DFF_P_  (.D(_00035_),
    .Q(\hash.CA1.w_i2[12] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[13]$_DFF_P_  (.D(_00036_),
    .Q(\hash.CA1.w_i2[13] ),
    .CLK(clknet_leaf_185_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[14]$_DFF_P_  (.D(_00037_),
    .Q(\hash.CA1.w_i2[14] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[15]$_DFF_P_  (.D(_00038_),
    .Q(\hash.CA1.w_i2[15] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[16]$_DFF_P_  (.D(_00039_),
    .Q(\hash.CA1.w_i2[16] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[17]$_DFF_P_  (.D(_00040_),
    .Q(\hash.CA1.w_i2[17] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[18]$_DFF_P_  (.D(_00041_),
    .Q(\hash.CA1.w_i2[18] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[19]$_DFF_P_  (.D(_00042_),
    .Q(\hash.CA1.w_i2[19] ),
    .CLK(clknet_leaf_234_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[1]$_DFF_P_  (.D(_00043_),
    .Q(\hash.CA1.w_i2[1] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[20]$_DFF_P_  (.D(_00044_),
    .Q(\hash.CA1.w_i2[20] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[21]$_DFF_P_  (.D(_00045_),
    .Q(\hash.CA1.w_i2[21] ),
    .CLK(clknet_leaf_233_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[22]$_DFF_P_  (.D(_00046_),
    .Q(\hash.CA1.w_i2[22] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[23]$_DFF_P_  (.D(_00047_),
    .Q(\hash.CA1.w_i2[23] ),
    .CLK(clknet_leaf_184_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[24]$_DFF_P_  (.D(_00048_),
    .Q(\hash.CA1.w_i2[24] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[25]$_DFF_P_  (.D(_00049_),
    .Q(\hash.CA1.w_i2[25] ),
    .CLK(clknet_leaf_231_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[26]$_DFF_P_  (.D(_00050_),
    .Q(\hash.CA1.w_i2[26] ),
    .CLK(clknet_leaf_181_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[27]$_DFF_P_  (.D(_00051_),
    .Q(\hash.CA1.w_i2[27] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[28]$_DFF_P_  (.D(_00052_),
    .Q(\hash.CA1.w_i2[28] ),
    .CLK(clknet_leaf_249_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[29]$_DFF_P_  (.D(_00053_),
    .Q(\hash.CA1.w_i2[29] ),
    .CLK(clknet_leaf_183_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[2]$_DFF_P_  (.D(_00054_),
    .Q(\hash.CA1.w_i2[2] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[30]$_DFF_P_  (.D(_00055_),
    .Q(\hash.CA1.w_i2[30] ),
    .CLK(clknet_leaf_182_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[31]$_DFF_P_  (.D(_00056_),
    .Q(\hash.CA1.w_i2[31] ),
    .CLK(clknet_leaf_236_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[3]$_DFF_P_  (.D(_00057_),
    .Q(\hash.CA1.w_i2[3] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[4]$_DFF_P_  (.D(_00058_),
    .Q(\hash.CA1.w_i2[4] ),
    .CLK(clknet_leaf_232_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[5]$_DFF_P_  (.D(_00059_),
    .Q(\hash.CA1.w_i2[5] ),
    .CLK(clknet_leaf_226_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[6]$_DFF_P_  (.D(_00060_),
    .Q(\hash.CA1.w_i2[6] ),
    .CLK(clknet_leaf_220_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[7]$_DFF_P_  (.D(_00061_),
    .Q(\hash.CA1.w_i2[7] ),
    .CLK(clknet_leaf_235_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[8]$_DFF_P_  (.D(_00062_),
    .Q(\hash.CA1.w_i2[8] ),
    .CLK(clknet_leaf_230_clk));
 sky130_fd_sc_hd__dfxtp_1 \w_value2[9]$_DFF_P_  (.D(_00063_),
    .Q(\hash.CA1.w_i2[9] ),
    .CLK(clknet_leaf_241_clk));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_212_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_213_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_214_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_215_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_216_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_217_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_218_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_219_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_220_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_221_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_222_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_223_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_224_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_225_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_226_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_227_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_228_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_229_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_230_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_231_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_232_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_233_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_234_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_235_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_236_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_237_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_238_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_239_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_240_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_241_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_242_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_243_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_244_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_245_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_246_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_247_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_248_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_249_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_250_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_251_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_252_6246 ();
 sky130_fd_sc_hd__buf_12 load_slew285 (.A(_09875_),
    .X(net285));
 sky130_fd_sc_hd__buf_12 load_slew286 (.A(net287),
    .X(net286));
 sky130_fd_sc_hd__buf_12 load_slew287 (.A(_09875_),
    .X(net287));
 sky130_fd_sc_hd__buf_12 load_slew288 (.A(net289),
    .X(net288));
 sky130_fd_sc_hd__buf_12 load_slew289 (.A(net290),
    .X(net289));
 sky130_fd_sc_hd__buf_12 load_slew290 (.A(_10373_),
    .X(net290));
 sky130_fd_sc_hd__buf_12 load_slew291 (.A(_10373_),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_4 wire292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__buf_12 load_slew293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_16 load_slew294 (.A(_09867_),
    .X(net294));
 sky130_fd_sc_hd__buf_12 load_slew295 (.A(_09867_),
    .X(net295));
 sky130_fd_sc_hd__buf_12 load_slew296 (.A(_00071_),
    .X(net296));
 sky130_fd_sc_hd__buf_12 max_cap297 (.A(_00071_),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_4 wire298 (.A(net300),
    .X(net298));
 sky130_fd_sc_hd__buf_12 load_slew299 (.A(net300),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_4 wire300 (.A(_00080_),
    .X(net300));
 sky130_fd_sc_hd__buf_12 load_slew301 (.A(net302),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_4 wire302 (.A(_00088_),
    .X(net302));
 sky130_fd_sc_hd__buf_12 max_cap303 (.A(net307),
    .X(net303));
 sky130_fd_sc_hd__buf_12 load_slew304 (.A(net306),
    .X(net304));
 sky130_fd_sc_hd__buf_12 load_slew305 (.A(net306),
    .X(net305));
 sky130_fd_sc_hd__buf_12 load_slew306 (.A(_00655_),
    .X(net306));
 sky130_fd_sc_hd__buf_12 load_slew307 (.A(_00655_),
    .X(net307));
 sky130_fd_sc_hd__buf_12 load_slew308 (.A(_00657_),
    .X(net308));
 sky130_fd_sc_hd__buf_12 load_slew309 (.A(net310),
    .X(net309));
 sky130_fd_sc_hd__buf_12 load_slew310 (.A(_00657_),
    .X(net310));
 sky130_fd_sc_hd__buf_12 load_slew311 (.A(_00657_),
    .X(net311));
 sky130_fd_sc_hd__buf_12 load_slew312 (.A(_00657_),
    .X(net312));
 sky130_fd_sc_hd__buf_12 max_cap313 (.A(net314),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_4 wire314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__buf_12 load_slew315 (.A(_10352_),
    .X(net315));
 sky130_fd_sc_hd__buf_12 load_slew316 (.A(net318),
    .X(net316));
 sky130_fd_sc_hd__buf_12 max_cap317 (.A(net318),
    .X(net317));
 sky130_fd_sc_hd__buf_12 max_cap318 (.A(_10352_),
    .X(net318));
 sky130_fd_sc_hd__buf_12 max_cap319 (.A(net320),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_4 wire320 (.A(_10348_),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_4 wire321 (.A(_10348_),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_4 wire322 (.A(net324),
    .X(net322));
 sky130_fd_sc_hd__buf_12 load_slew323 (.A(net324),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_4 wire324 (.A(net325),
    .X(net324));
 sky130_fd_sc_hd__buf_12 load_slew325 (.A(_10348_),
    .X(net325));
 sky130_fd_sc_hd__buf_12 load_slew326 (.A(net328),
    .X(net326));
 sky130_fd_sc_hd__buf_12 max_cap327 (.A(net328),
    .X(net327));
 sky130_fd_sc_hd__buf_12 load_slew328 (.A(_09857_),
    .X(net328));
 sky130_fd_sc_hd__buf_12 load_slew329 (.A(_09857_),
    .X(net329));
 sky130_fd_sc_hd__buf_12 load_slew330 (.A(net331),
    .X(net330));
 sky130_fd_sc_hd__buf_12 max_cap331 (.A(_09857_),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_4 wire332 (.A(_09854_),
    .X(net332));
 sky130_fd_sc_hd__buf_12 load_slew333 (.A(net334),
    .X(net333));
 sky130_fd_sc_hd__buf_12 max_cap334 (.A(net337),
    .X(net334));
 sky130_fd_sc_hd__buf_12 max_cap335 (.A(net336),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_4 wire336 (.A(net338),
    .X(net336));
 sky130_fd_sc_hd__buf_12 load_slew337 (.A(net338),
    .X(net337));
 sky130_fd_sc_hd__buf_12 load_slew338 (.A(_09854_),
    .X(net338));
 sky130_fd_sc_hd__buf_12 load_slew339 (.A(_04797_),
    .X(net339));
 sky130_fd_sc_hd__buf_12 load_slew340 (.A(net341),
    .X(net340));
 sky130_fd_sc_hd__buf_12 load_slew341 (.A(net346),
    .X(net341));
 sky130_fd_sc_hd__buf_12 load_slew342 (.A(net345),
    .X(net342));
 sky130_fd_sc_hd__buf_12 load_slew343 (.A(net344),
    .X(net343));
 sky130_fd_sc_hd__buf_12 load_slew344 (.A(net345),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_1 load_slew345 (.A(net534),
    .X(net345));
 sky130_fd_sc_hd__buf_12 max_cap346 (.A(\hash.reset ),
    .X(net346));
 sky130_fd_sc_hd__buf_12 load_slew347 (.A(net349),
    .X(net347));
 sky130_fd_sc_hd__buf_12 load_slew348 (.A(reset_hash),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_1 load_slew349 (.A(reset_hash),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_4 wire350 (.A(net351),
    .X(net350));
 sky130_fd_sc_hd__buf_12 load_slew351 (.A(net355),
    .X(net351));
 sky130_fd_sc_hd__buf_12 load_slew352 (.A(net355),
    .X(net352));
 sky130_fd_sc_hd__buf_12 load_slew353 (.A(net354),
    .X(net353));
 sky130_fd_sc_hd__buf_12 load_slew354 (.A(net356),
    .X(net354));
 sky130_fd_sc_hd__buf_12 load_slew355 (.A(net356),
    .X(net355));
 sky130_fd_sc_hd__buf_12 load_slew356 (.A(done),
    .X(net356));
 sky130_fd_sc_hd__buf_12 load_slew357 (.A(net364),
    .X(net357));
 sky130_fd_sc_hd__buf_12 load_slew358 (.A(net362),
    .X(net358));
 sky130_fd_sc_hd__buf_12 load_slew359 (.A(net362),
    .X(net359));
 sky130_fd_sc_hd__buf_12 load_slew360 (.A(net362),
    .X(net360));
 sky130_fd_sc_hd__buf_12 load_slew361 (.A(net363),
    .X(net361));
 sky130_fd_sc_hd__buf_12 load_slew362 (.A(net363),
    .X(net362));
 sky130_fd_sc_hd__buf_12 max_cap363 (.A(net364),
    .X(net363));
 sky130_fd_sc_hd__buf_12 load_slew364 (.A(\count_hash2[1] ),
    .X(net364));
 sky130_fd_sc_hd__buf_12 load_slew365 (.A(net366),
    .X(net365));
 sky130_fd_sc_hd__buf_12 load_slew366 (.A(net370),
    .X(net366));
 sky130_fd_sc_hd__buf_12 load_slew367 (.A(net368),
    .X(net367));
 sky130_fd_sc_hd__buf_12 load_slew368 (.A(net370),
    .X(net368));
 sky130_fd_sc_hd__buf_12 load_slew369 (.A(net372),
    .X(net369));
 sky130_fd_sc_hd__buf_12 load_slew370 (.A(net372),
    .X(net370));
 sky130_fd_sc_hd__buf_12 load_slew371 (.A(\count_hash1[1] ),
    .X(net371));
 sky130_fd_sc_hd__buf_12 load_slew372 (.A(\count_hash1[1] ),
    .X(net372));
 sky130_fd_sc_hd__buf_12 load_slew373 (.A(net374),
    .X(net373));
 sky130_fd_sc_hd__buf_12 load_slew374 (.A(\count7_2[5] ),
    .X(net374));
 sky130_fd_sc_hd__buf_12 load_slew375 (.A(net376),
    .X(net375));
 sky130_fd_sc_hd__buf_12 load_slew376 (.A(\count7_2[4] ),
    .X(net376));
 sky130_fd_sc_hd__buf_12 load_slew377 (.A(net379),
    .X(net377));
 sky130_fd_sc_hd__buf_12 load_slew378 (.A(net379),
    .X(net378));
 sky130_fd_sc_hd__buf_12 load_slew379 (.A(\count7_2[3] ),
    .X(net379));
 sky130_fd_sc_hd__buf_12 load_slew380 (.A(net387),
    .X(net380));
 sky130_fd_sc_hd__buf_12 load_slew381 (.A(net382),
    .X(net381));
 sky130_fd_sc_hd__buf_12 load_slew382 (.A(net383),
    .X(net382));
 sky130_fd_sc_hd__buf_12 load_slew383 (.A(net385),
    .X(net383));
 sky130_fd_sc_hd__buf_12 max_cap384 (.A(net385),
    .X(net384));
 sky130_fd_sc_hd__buf_12 max_cap385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__buf_12 load_slew386 (.A(\count7_2[2] ),
    .X(net386));
 sky130_fd_sc_hd__buf_12 load_slew387 (.A(\count7_2[2] ),
    .X(net387));
 sky130_fd_sc_hd__buf_12 load_slew388 (.A(\count7_2[1] ),
    .X(net388));
 sky130_fd_sc_hd__buf_12 load_slew389 (.A(net390),
    .X(net389));
 sky130_fd_sc_hd__buf_12 load_slew390 (.A(net392),
    .X(net390));
 sky130_fd_sc_hd__buf_12 load_slew391 (.A(net392),
    .X(net391));
 sky130_fd_sc_hd__buf_12 load_slew392 (.A(net393),
    .X(net392));
 sky130_fd_sc_hd__buf_12 load_slew393 (.A(\count7_2[1] ),
    .X(net393));
 sky130_fd_sc_hd__buf_12 load_slew394 (.A(net395),
    .X(net394));
 sky130_fd_sc_hd__buf_12 load_slew395 (.A(\count7_1[5] ),
    .X(net395));
 sky130_fd_sc_hd__buf_12 load_slew396 (.A(net536),
    .X(net396));
 sky130_fd_sc_hd__buf_12 load_slew397 (.A(net536),
    .X(net397));
 sky130_fd_sc_hd__buf_12 load_slew398 (.A(net537),
    .X(net398));
 sky130_fd_sc_hd__buf_12 load_slew399 (.A(net537),
    .X(net399));
 sky130_fd_sc_hd__buf_12 load_slew400 (.A(\count7_1[3] ),
    .X(net400));
 sky130_fd_sc_hd__buf_12 load_slew401 (.A(net405),
    .X(net401));
 sky130_fd_sc_hd__buf_12 load_slew402 (.A(net404),
    .X(net402));
 sky130_fd_sc_hd__buf_12 load_slew403 (.A(net404),
    .X(net403));
 sky130_fd_sc_hd__buf_12 load_slew404 (.A(net406),
    .X(net404));
 sky130_fd_sc_hd__buf_12 load_slew405 (.A(net406),
    .X(net405));
 sky130_fd_sc_hd__buf_12 load_slew406 (.A(\count7_1[2] ),
    .X(net406));
 sky130_fd_sc_hd__buf_12 load_slew407 (.A(\count7_1[2] ),
    .X(net407));
 sky130_fd_sc_hd__buf_12 load_slew408 (.A(net409),
    .X(net408));
 sky130_fd_sc_hd__buf_12 load_slew409 (.A(\count7_1[1] ),
    .X(net409));
 sky130_fd_sc_hd__buf_12 load_slew410 (.A(net411),
    .X(net410));
 sky130_fd_sc_hd__buf_12 load_slew411 (.A(net412),
    .X(net411));
 sky130_fd_sc_hd__buf_12 load_slew412 (.A(\count7_1[1] ),
    .X(net412));
 sky130_fd_sc_hd__buf_12 max_cap413 (.A(\count2_2[5] ),
    .X(net413));
 sky130_fd_sc_hd__buf_12 load_slew414 (.A(net540),
    .X(net414));
 sky130_fd_sc_hd__buf_12 load_slew415 (.A(\count2_2[4] ),
    .X(net415));
 sky130_fd_sc_hd__buf_12 load_slew416 (.A(net417),
    .X(net416));
 sky130_fd_sc_hd__buf_12 load_slew417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__buf_12 load_slew418 (.A(\count2_2[3] ),
    .X(net418));
 sky130_fd_sc_hd__buf_12 load_slew419 (.A(net421),
    .X(net419));
 sky130_fd_sc_hd__buf_12 load_slew420 (.A(net423),
    .X(net420));
 sky130_fd_sc_hd__buf_12 load_slew421 (.A(net423),
    .X(net421));
 sky130_fd_sc_hd__buf_12 load_slew422 (.A(net424),
    .X(net422));
 sky130_fd_sc_hd__buf_12 max_cap423 (.A(net424),
    .X(net423));
 sky130_fd_sc_hd__buf_12 load_slew424 (.A(net541),
    .X(net424));
 sky130_fd_sc_hd__buf_12 load_slew425 (.A(\count2_2[2] ),
    .X(net425));
 sky130_fd_sc_hd__buf_12 load_slew426 (.A(net428),
    .X(net426));
 sky130_fd_sc_hd__buf_12 load_slew427 (.A(net428),
    .X(net427));
 sky130_fd_sc_hd__buf_12 load_slew428 (.A(net429),
    .X(net428));
 sky130_fd_sc_hd__buf_12 load_slew429 (.A(net430),
    .X(net429));
 sky130_fd_sc_hd__buf_12 load_slew430 (.A(net431),
    .X(net430));
 sky130_fd_sc_hd__buf_12 load_slew431 (.A(\count2_2[1] ),
    .X(net431));
 sky130_fd_sc_hd__buf_12 load_slew432 (.A(net433),
    .X(net432));
 sky130_fd_sc_hd__buf_12 load_slew433 (.A(\count2_1[5] ),
    .X(net433));
 sky130_fd_sc_hd__buf_12 load_slew434 (.A(net435),
    .X(net434));
 sky130_fd_sc_hd__buf_12 load_slew435 (.A(\count2_1[4] ),
    .X(net435));
 sky130_fd_sc_hd__buf_12 load_slew436 (.A(net438),
    .X(net436));
 sky130_fd_sc_hd__buf_12 load_slew437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__buf_12 load_slew438 (.A(\count2_1[3] ),
    .X(net438));
 sky130_fd_sc_hd__buf_12 load_slew439 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__buf_12 load_slew440 (.A(net441),
    .X(net440));
 sky130_fd_sc_hd__buf_12 load_slew441 (.A(net443),
    .X(net441));
 sky130_fd_sc_hd__buf_12 load_slew442 (.A(net443),
    .X(net442));
 sky130_fd_sc_hd__buf_12 max_cap443 (.A(net445),
    .X(net443));
 sky130_fd_sc_hd__buf_12 load_slew444 (.A(net446),
    .X(net444));
 sky130_fd_sc_hd__buf_12 max_cap445 (.A(net446),
    .X(net445));
 sky130_fd_sc_hd__buf_12 load_slew446 (.A(\count2_1[2] ),
    .X(net446));
 sky130_fd_sc_hd__buf_12 load_slew447 (.A(\count2_1[1] ),
    .X(net447));
 sky130_fd_sc_hd__buf_12 load_slew448 (.A(net449),
    .X(net448));
 sky130_fd_sc_hd__buf_12 load_slew449 (.A(net451),
    .X(net449));
 sky130_fd_sc_hd__buf_12 load_slew450 (.A(net451),
    .X(net450));
 sky130_fd_sc_hd__buf_12 load_slew451 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__buf_12 load_slew452 (.A(net1093),
    .X(net452));
 sky130_fd_sc_hd__buf_12 load_slew453 (.A(net542),
    .X(net453));
 sky130_fd_sc_hd__buf_12 load_slew454 (.A(net543),
    .X(net454));
 sky130_fd_sc_hd__buf_12 load_slew455 (.A(net543),
    .X(net455));
 sky130_fd_sc_hd__buf_12 load_slew456 (.A(\count16_2[3] ),
    .X(net456));
 sky130_fd_sc_hd__buf_12 load_slew457 (.A(\count16_2[3] ),
    .X(net457));
 sky130_fd_sc_hd__buf_12 load_slew458 (.A(\count16_2[3] ),
    .X(net458));
 sky130_fd_sc_hd__buf_12 load_slew459 (.A(net460),
    .X(net459));
 sky130_fd_sc_hd__buf_12 load_slew460 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__buf_12 load_slew461 (.A(net462),
    .X(net461));
 sky130_fd_sc_hd__buf_12 load_slew462 (.A(net466),
    .X(net462));
 sky130_fd_sc_hd__buf_12 load_slew463 (.A(net465),
    .X(net463));
 sky130_fd_sc_hd__buf_12 load_slew464 (.A(net465),
    .X(net464));
 sky130_fd_sc_hd__buf_12 load_slew465 (.A(\count16_2[2] ),
    .X(net465));
 sky130_fd_sc_hd__buf_12 load_slew466 (.A(\count16_2[2] ),
    .X(net466));
 sky130_fd_sc_hd__buf_12 load_slew467 (.A(net469),
    .X(net467));
 sky130_fd_sc_hd__buf_12 load_slew468 (.A(net469),
    .X(net468));
 sky130_fd_sc_hd__buf_12 load_slew469 (.A(net470),
    .X(net469));
 sky130_fd_sc_hd__buf_12 load_slew470 (.A(net471),
    .X(net470));
 sky130_fd_sc_hd__buf_12 load_slew471 (.A(\count16_2[1] ),
    .X(net471));
 sky130_fd_sc_hd__buf_12 load_slew472 (.A(net473),
    .X(net472));
 sky130_fd_sc_hd__buf_12 load_slew473 (.A(net545),
    .X(net473));
 sky130_fd_sc_hd__buf_12 load_slew474 (.A(\count16_1[4] ),
    .X(net474));
 sky130_fd_sc_hd__buf_12 load_slew475 (.A(\count16_1[4] ),
    .X(net475));
 sky130_fd_sc_hd__buf_12 load_slew476 (.A(net546),
    .X(net476));
 sky130_fd_sc_hd__buf_12 load_slew477 (.A(\count16_1[3] ),
    .X(net477));
 sky130_fd_sc_hd__buf_12 load_slew478 (.A(net485),
    .X(net478));
 sky130_fd_sc_hd__buf_12 load_slew479 (.A(net480),
    .X(net479));
 sky130_fd_sc_hd__buf_12 load_slew480 (.A(net481),
    .X(net480));
 sky130_fd_sc_hd__buf_12 load_slew481 (.A(net482),
    .X(net481));
 sky130_fd_sc_hd__buf_12 load_slew482 (.A(net483),
    .X(net482));
 sky130_fd_sc_hd__buf_12 load_slew483 (.A(\count16_1[2] ),
    .X(net483));
 sky130_fd_sc_hd__buf_12 load_slew484 (.A(\count16_1[2] ),
    .X(net484));
 sky130_fd_sc_hd__buf_12 load_slew485 (.A(\count16_1[2] ),
    .X(net485));
 sky130_fd_sc_hd__buf_12 load_slew486 (.A(\count16_1[1] ),
    .X(net486));
 sky130_fd_sc_hd__buf_12 load_slew487 (.A(net488),
    .X(net487));
 sky130_fd_sc_hd__buf_12 load_slew488 (.A(net491),
    .X(net488));
 sky130_fd_sc_hd__buf_12 load_slew489 (.A(net490),
    .X(net489));
 sky130_fd_sc_hd__buf_12 max_cap490 (.A(net491),
    .X(net490));
 sky130_fd_sc_hd__buf_12 load_slew491 (.A(\count16_1[1] ),
    .X(net491));
 sky130_fd_sc_hd__buf_12 load_slew492 (.A(net493),
    .X(net492));
 sky130_fd_sc_hd__buf_12 load_slew493 (.A(\count15_2[5] ),
    .X(net493));
 sky130_fd_sc_hd__buf_12 load_slew494 (.A(net547),
    .X(net494));
 sky130_fd_sc_hd__buf_12 load_slew495 (.A(\count15_2[4] ),
    .X(net495));
 sky130_fd_sc_hd__buf_12 load_slew496 (.A(\count15_2[3] ),
    .X(net496));
 sky130_fd_sc_hd__buf_12 load_slew497 (.A(net548),
    .X(net497));
 sky130_fd_sc_hd__buf_12 load_slew498 (.A(net499),
    .X(net498));
 sky130_fd_sc_hd__buf_12 load_slew499 (.A(\count15_2[2] ),
    .X(net499));
 sky130_fd_sc_hd__buf_12 load_slew500 (.A(net501),
    .X(net500));
 sky130_fd_sc_hd__buf_12 load_slew501 (.A(net502),
    .X(net501));
 sky130_fd_sc_hd__buf_12 load_slew502 (.A(net504),
    .X(net502));
 sky130_fd_sc_hd__buf_12 load_slew503 (.A(net504),
    .X(net503));
 sky130_fd_sc_hd__buf_16 load_slew504 (.A(net505),
    .X(net504));
 sky130_fd_sc_hd__buf_12 load_slew505 (.A(\count15_2[2] ),
    .X(net505));
 sky130_fd_sc_hd__buf_12 load_slew506 (.A(\count15_2[1] ),
    .X(net506));
 sky130_fd_sc_hd__buf_12 load_slew507 (.A(net508),
    .X(net507));
 sky130_fd_sc_hd__buf_12 load_slew508 (.A(net510),
    .X(net508));
 sky130_fd_sc_hd__buf_12 load_slew509 (.A(net510),
    .X(net509));
 sky130_fd_sc_hd__buf_12 load_slew510 (.A(net511),
    .X(net510));
 sky130_fd_sc_hd__buf_12 load_slew511 (.A(\count15_2[1] ),
    .X(net511));
 sky130_fd_sc_hd__buf_12 load_slew512 (.A(net513),
    .X(net512));
 sky130_fd_sc_hd__buf_12 load_slew513 (.A(\count15_1[5] ),
    .X(net513));
 sky130_fd_sc_hd__buf_12 load_slew514 (.A(net549),
    .X(net514));
 sky130_fd_sc_hd__buf_12 load_slew515 (.A(\count15_1[4] ),
    .X(net515));
 sky130_fd_sc_hd__buf_12 load_slew516 (.A(net518),
    .X(net516));
 sky130_fd_sc_hd__buf_12 load_slew517 (.A(\count15_1[3] ),
    .X(net517));
 sky130_fd_sc_hd__buf_12 load_slew518 (.A(\count15_1[3] ),
    .X(net518));
 sky130_fd_sc_hd__buf_12 load_slew519 (.A(net523),
    .X(net519));
 sky130_fd_sc_hd__buf_12 load_slew520 (.A(net521),
    .X(net520));
 sky130_fd_sc_hd__buf_12 load_slew521 (.A(net522),
    .X(net521));
 sky130_fd_sc_hd__buf_12 load_slew522 (.A(net523),
    .X(net522));
 sky130_fd_sc_hd__buf_12 load_slew523 (.A(\count15_1[2] ),
    .X(net523));
 sky130_fd_sc_hd__buf_12 load_slew524 (.A(net525),
    .X(net524));
 sky130_fd_sc_hd__buf_12 load_slew525 (.A(net526),
    .X(net525));
 sky130_fd_sc_hd__buf_12 load_slew526 (.A(net527),
    .X(net526));
 sky130_fd_sc_hd__buf_12 load_slew527 (.A(\count15_1[2] ),
    .X(net527));
 sky130_fd_sc_hd__buf_12 load_slew528 (.A(net532),
    .X(net528));
 sky130_fd_sc_hd__buf_12 load_slew529 (.A(net531),
    .X(net529));
 sky130_fd_sc_hd__buf_12 load_slew530 (.A(net531),
    .X(net530));
 sky130_fd_sc_hd__buf_12 load_slew531 (.A(net532),
    .X(net531));
 sky130_fd_sc_hd__buf_12 load_slew532 (.A(\count15_1[1] ),
    .X(net532));
 sky130_fd_sc_hd__buf_12 load_slew533 (.A(_08591_),
    .X(net533));
 sky130_fd_sc_hd__buf_12 load_slew534 (.A(\hash.reset ),
    .X(net534));
 sky130_fd_sc_hd__buf_12 load_slew535 (.A(\count7_2[4] ),
    .X(net535));
 sky130_fd_sc_hd__buf_12 load_slew536 (.A(\count7_1[4] ),
    .X(net536));
 sky130_fd_sc_hd__buf_12 load_slew537 (.A(\count7_1[3] ),
    .X(net537));
 sky130_fd_sc_hd__buf_12 load_slew538 (.A(\count7_1[2] ),
    .X(net538));
 sky130_fd_sc_hd__buf_12 load_slew539 (.A(\count2_2[5] ),
    .X(net539));
 sky130_fd_sc_hd__buf_12 load_slew540 (.A(\count2_2[4] ),
    .X(net540));
 sky130_fd_sc_hd__buf_12 load_slew541 (.A(\count2_2[2] ),
    .X(net541));
 sky130_fd_sc_hd__buf_12 load_slew542 (.A(\count16_2[5] ),
    .X(net542));
 sky130_fd_sc_hd__buf_12 load_slew543 (.A(\count16_2[4] ),
    .X(net543));
 sky130_fd_sc_hd__buf_12 load_slew544 (.A(\count16_2[1] ),
    .X(net544));
 sky130_fd_sc_hd__buf_12 load_slew545 (.A(\count16_1[5] ),
    .X(net545));
 sky130_fd_sc_hd__buf_12 load_slew546 (.A(\count16_1[3] ),
    .X(net546));
 sky130_fd_sc_hd__buf_12 load_slew547 (.A(\count15_2[4] ),
    .X(net547));
 sky130_fd_sc_hd__buf_12 load_slew548 (.A(\count15_2[3] ),
    .X(net548));
 sky130_fd_sc_hd__buf_12 load_slew549 (.A(\count15_1[4] ),
    .X(net549));
 sky130_fd_sc_hd__buf_12 load_slew550 (.A(\count15_1[1] ),
    .X(net550));
 sky130_fd_sc_hd__buf_12 load_slew551 (.A(_09784_),
    .X(net551));
 sky130_fd_sc_hd__buf_1 input1 (.A(message[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(message[100]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(message[101]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(message[102]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(message[103]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(message[104]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(message[105]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(message[106]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(message[107]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(message[108]),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(message[109]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(message[10]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(message[110]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(message[111]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(message[112]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(message[113]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(message[114]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(message[115]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(message[116]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input20 (.A(message[117]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(message[118]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(message[119]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(message[11]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(message[120]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(message[121]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(message[122]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(message[123]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(message[124]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(message[125]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(message[126]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(message[127]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(message[128]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(message[129]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(message[12]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(message[130]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(message[131]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(message[132]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(message[133]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(message[134]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input40 (.A(message[135]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(message[136]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(message[137]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(message[138]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(message[139]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(message[13]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(message[140]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(message[141]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(message[142]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(message[143]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input50 (.A(message[144]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(message[145]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(message[146]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(message[147]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(message[148]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(message[149]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(message[14]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(message[150]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(message[151]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(message[152]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input60 (.A(message[153]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(message[154]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(message[155]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(message[156]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(message[157]),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(message[158]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(message[159]),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input67 (.A(message[15]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(message[160]),
    .X(net68));
 sky130_fd_sc_hd__buf_1 input69 (.A(message[161]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input70 (.A(message[162]),
    .X(net70));
 sky130_fd_sc_hd__buf_1 input71 (.A(message[163]),
    .X(net71));
 sky130_fd_sc_hd__buf_1 input72 (.A(message[164]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(message[165]),
    .X(net73));
 sky130_fd_sc_hd__buf_1 input74 (.A(message[166]),
    .X(net74));
 sky130_fd_sc_hd__buf_1 input75 (.A(message[167]),
    .X(net75));
 sky130_fd_sc_hd__buf_1 input76 (.A(message[168]),
    .X(net76));
 sky130_fd_sc_hd__buf_1 input77 (.A(message[169]),
    .X(net77));
 sky130_fd_sc_hd__buf_1 input78 (.A(message[16]),
    .X(net78));
 sky130_fd_sc_hd__buf_1 input79 (.A(message[170]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input80 (.A(message[171]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input81 (.A(message[172]),
    .X(net81));
 sky130_fd_sc_hd__buf_1 input82 (.A(message[173]),
    .X(net82));
 sky130_fd_sc_hd__buf_1 input83 (.A(message[174]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 input84 (.A(message[175]),
    .X(net84));
 sky130_fd_sc_hd__buf_1 input85 (.A(message[176]),
    .X(net85));
 sky130_fd_sc_hd__buf_1 input86 (.A(message[177]),
    .X(net86));
 sky130_fd_sc_hd__buf_1 input87 (.A(message[178]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 input88 (.A(message[179]),
    .X(net88));
 sky130_fd_sc_hd__buf_1 input89 (.A(message[17]),
    .X(net89));
 sky130_fd_sc_hd__buf_1 input90 (.A(message[180]),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input91 (.A(message[181]),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input92 (.A(message[182]),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input93 (.A(message[183]),
    .X(net93));
 sky130_fd_sc_hd__buf_1 input94 (.A(message[184]),
    .X(net94));
 sky130_fd_sc_hd__buf_1 input95 (.A(message[185]),
    .X(net95));
 sky130_fd_sc_hd__buf_1 input96 (.A(message[186]),
    .X(net96));
 sky130_fd_sc_hd__buf_1 input97 (.A(message[187]),
    .X(net97));
 sky130_fd_sc_hd__buf_1 input98 (.A(message[188]),
    .X(net98));
 sky130_fd_sc_hd__buf_1 input99 (.A(message[189]),
    .X(net99));
 sky130_fd_sc_hd__buf_1 input100 (.A(message[18]),
    .X(net100));
 sky130_fd_sc_hd__buf_1 input101 (.A(message[190]),
    .X(net101));
 sky130_fd_sc_hd__buf_1 input102 (.A(message[191]),
    .X(net102));
 sky130_fd_sc_hd__buf_1 input103 (.A(message[192]),
    .X(net103));
 sky130_fd_sc_hd__buf_1 input104 (.A(message[193]),
    .X(net104));
 sky130_fd_sc_hd__buf_1 input105 (.A(message[194]),
    .X(net105));
 sky130_fd_sc_hd__buf_1 input106 (.A(message[195]),
    .X(net106));
 sky130_fd_sc_hd__buf_1 input107 (.A(message[196]),
    .X(net107));
 sky130_fd_sc_hd__buf_1 input108 (.A(message[197]),
    .X(net108));
 sky130_fd_sc_hd__buf_1 input109 (.A(message[198]),
    .X(net109));
 sky130_fd_sc_hd__buf_1 input110 (.A(message[199]),
    .X(net110));
 sky130_fd_sc_hd__buf_1 input111 (.A(message[19]),
    .X(net111));
 sky130_fd_sc_hd__buf_1 input112 (.A(message[1]),
    .X(net112));
 sky130_fd_sc_hd__buf_1 input113 (.A(message[200]),
    .X(net113));
 sky130_fd_sc_hd__buf_1 input114 (.A(message[201]),
    .X(net114));
 sky130_fd_sc_hd__buf_1 input115 (.A(message[202]),
    .X(net115));
 sky130_fd_sc_hd__buf_1 input116 (.A(message[203]),
    .X(net116));
 sky130_fd_sc_hd__buf_1 input117 (.A(message[204]),
    .X(net117));
 sky130_fd_sc_hd__buf_1 input118 (.A(message[205]),
    .X(net118));
 sky130_fd_sc_hd__buf_1 input119 (.A(message[206]),
    .X(net119));
 sky130_fd_sc_hd__buf_1 input120 (.A(message[207]),
    .X(net120));
 sky130_fd_sc_hd__buf_1 input121 (.A(message[208]),
    .X(net121));
 sky130_fd_sc_hd__buf_1 input122 (.A(message[209]),
    .X(net122));
 sky130_fd_sc_hd__buf_1 input123 (.A(message[20]),
    .X(net123));
 sky130_fd_sc_hd__buf_1 input124 (.A(message[210]),
    .X(net124));
 sky130_fd_sc_hd__buf_1 input125 (.A(message[211]),
    .X(net125));
 sky130_fd_sc_hd__buf_1 input126 (.A(message[212]),
    .X(net126));
 sky130_fd_sc_hd__buf_1 input127 (.A(message[213]),
    .X(net127));
 sky130_fd_sc_hd__buf_1 input128 (.A(message[214]),
    .X(net128));
 sky130_fd_sc_hd__buf_1 input129 (.A(message[215]),
    .X(net129));
 sky130_fd_sc_hd__buf_1 input130 (.A(message[216]),
    .X(net130));
 sky130_fd_sc_hd__buf_1 input131 (.A(message[217]),
    .X(net131));
 sky130_fd_sc_hd__buf_1 input132 (.A(message[218]),
    .X(net132));
 sky130_fd_sc_hd__buf_1 input133 (.A(message[219]),
    .X(net133));
 sky130_fd_sc_hd__buf_1 input134 (.A(message[21]),
    .X(net134));
 sky130_fd_sc_hd__buf_1 input135 (.A(message[220]),
    .X(net135));
 sky130_fd_sc_hd__buf_1 input136 (.A(message[221]),
    .X(net136));
 sky130_fd_sc_hd__buf_1 input137 (.A(message[222]),
    .X(net137));
 sky130_fd_sc_hd__buf_1 input138 (.A(message[223]),
    .X(net138));
 sky130_fd_sc_hd__buf_1 input139 (.A(message[224]),
    .X(net139));
 sky130_fd_sc_hd__buf_1 input140 (.A(message[225]),
    .X(net140));
 sky130_fd_sc_hd__buf_1 input141 (.A(message[226]),
    .X(net141));
 sky130_fd_sc_hd__buf_1 input142 (.A(message[227]),
    .X(net142));
 sky130_fd_sc_hd__buf_1 input143 (.A(message[228]),
    .X(net143));
 sky130_fd_sc_hd__buf_1 input144 (.A(message[229]),
    .X(net144));
 sky130_fd_sc_hd__buf_1 input145 (.A(message[22]),
    .X(net145));
 sky130_fd_sc_hd__buf_1 input146 (.A(message[230]),
    .X(net146));
 sky130_fd_sc_hd__buf_1 input147 (.A(message[231]),
    .X(net147));
 sky130_fd_sc_hd__buf_1 input148 (.A(message[232]),
    .X(net148));
 sky130_fd_sc_hd__buf_1 input149 (.A(message[233]),
    .X(net149));
 sky130_fd_sc_hd__buf_1 input150 (.A(message[234]),
    .X(net150));
 sky130_fd_sc_hd__buf_1 input151 (.A(message[235]),
    .X(net151));
 sky130_fd_sc_hd__buf_1 input152 (.A(message[236]),
    .X(net152));
 sky130_fd_sc_hd__buf_1 input153 (.A(message[237]),
    .X(net153));
 sky130_fd_sc_hd__buf_1 input154 (.A(message[238]),
    .X(net154));
 sky130_fd_sc_hd__buf_1 input155 (.A(message[239]),
    .X(net155));
 sky130_fd_sc_hd__buf_1 input156 (.A(message[23]),
    .X(net156));
 sky130_fd_sc_hd__buf_1 input157 (.A(message[240]),
    .X(net157));
 sky130_fd_sc_hd__buf_1 input158 (.A(message[241]),
    .X(net158));
 sky130_fd_sc_hd__buf_1 input159 (.A(message[242]),
    .X(net159));
 sky130_fd_sc_hd__buf_1 input160 (.A(message[243]),
    .X(net160));
 sky130_fd_sc_hd__buf_1 input161 (.A(message[244]),
    .X(net161));
 sky130_fd_sc_hd__buf_1 input162 (.A(message[245]),
    .X(net162));
 sky130_fd_sc_hd__buf_1 input163 (.A(message[246]),
    .X(net163));
 sky130_fd_sc_hd__buf_1 input164 (.A(message[247]),
    .X(net164));
 sky130_fd_sc_hd__buf_1 input165 (.A(message[248]),
    .X(net165));
 sky130_fd_sc_hd__buf_1 input166 (.A(message[249]),
    .X(net166));
 sky130_fd_sc_hd__buf_1 input167 (.A(message[24]),
    .X(net167));
 sky130_fd_sc_hd__buf_1 input168 (.A(message[250]),
    .X(net168));
 sky130_fd_sc_hd__buf_1 input169 (.A(message[251]),
    .X(net169));
 sky130_fd_sc_hd__buf_1 input170 (.A(message[252]),
    .X(net170));
 sky130_fd_sc_hd__buf_1 input171 (.A(message[253]),
    .X(net171));
 sky130_fd_sc_hd__buf_1 input172 (.A(message[254]),
    .X(net172));
 sky130_fd_sc_hd__buf_1 input173 (.A(message[255]),
    .X(net173));
 sky130_fd_sc_hd__buf_1 input174 (.A(message[256]),
    .X(net174));
 sky130_fd_sc_hd__buf_1 input175 (.A(message[257]),
    .X(net175));
 sky130_fd_sc_hd__buf_1 input176 (.A(message[258]),
    .X(net176));
 sky130_fd_sc_hd__buf_1 input177 (.A(message[259]),
    .X(net177));
 sky130_fd_sc_hd__buf_1 input178 (.A(message[25]),
    .X(net178));
 sky130_fd_sc_hd__buf_1 input179 (.A(message[260]),
    .X(net179));
 sky130_fd_sc_hd__buf_1 input180 (.A(message[261]),
    .X(net180));
 sky130_fd_sc_hd__buf_1 input181 (.A(message[262]),
    .X(net181));
 sky130_fd_sc_hd__buf_1 input182 (.A(message[263]),
    .X(net182));
 sky130_fd_sc_hd__buf_1 input183 (.A(message[264]),
    .X(net183));
 sky130_fd_sc_hd__buf_1 input184 (.A(message[265]),
    .X(net184));
 sky130_fd_sc_hd__buf_1 input185 (.A(message[266]),
    .X(net185));
 sky130_fd_sc_hd__buf_1 input186 (.A(message[267]),
    .X(net186));
 sky130_fd_sc_hd__buf_1 input187 (.A(message[268]),
    .X(net187));
 sky130_fd_sc_hd__buf_1 input188 (.A(message[269]),
    .X(net188));
 sky130_fd_sc_hd__buf_1 input189 (.A(message[26]),
    .X(net189));
 sky130_fd_sc_hd__buf_1 input190 (.A(message[270]),
    .X(net190));
 sky130_fd_sc_hd__buf_1 input191 (.A(message[271]),
    .X(net191));
 sky130_fd_sc_hd__buf_1 input192 (.A(message[272]),
    .X(net192));
 sky130_fd_sc_hd__buf_1 input193 (.A(message[273]),
    .X(net193));
 sky130_fd_sc_hd__buf_1 input194 (.A(message[274]),
    .X(net194));
 sky130_fd_sc_hd__buf_1 input195 (.A(message[275]),
    .X(net195));
 sky130_fd_sc_hd__buf_1 input196 (.A(message[276]),
    .X(net196));
 sky130_fd_sc_hd__buf_1 input197 (.A(message[277]),
    .X(net197));
 sky130_fd_sc_hd__buf_1 input198 (.A(message[278]),
    .X(net198));
 sky130_fd_sc_hd__buf_1 input199 (.A(message[279]),
    .X(net199));
 sky130_fd_sc_hd__buf_1 input200 (.A(message[27]),
    .X(net200));
 sky130_fd_sc_hd__buf_1 input201 (.A(message[280]),
    .X(net201));
 sky130_fd_sc_hd__buf_1 input202 (.A(message[281]),
    .X(net202));
 sky130_fd_sc_hd__buf_1 input203 (.A(message[282]),
    .X(net203));
 sky130_fd_sc_hd__buf_1 input204 (.A(message[283]),
    .X(net204));
 sky130_fd_sc_hd__buf_1 input205 (.A(message[284]),
    .X(net205));
 sky130_fd_sc_hd__buf_1 input206 (.A(message[285]),
    .X(net206));
 sky130_fd_sc_hd__buf_1 input207 (.A(message[286]),
    .X(net207));
 sky130_fd_sc_hd__buf_1 input208 (.A(message[287]),
    .X(net208));
 sky130_fd_sc_hd__buf_1 input209 (.A(message[288]),
    .X(net209));
 sky130_fd_sc_hd__buf_1 input210 (.A(message[289]),
    .X(net210));
 sky130_fd_sc_hd__buf_1 input211 (.A(message[28]),
    .X(net211));
 sky130_fd_sc_hd__buf_1 input212 (.A(message[290]),
    .X(net212));
 sky130_fd_sc_hd__buf_1 input213 (.A(message[291]),
    .X(net213));
 sky130_fd_sc_hd__buf_1 input214 (.A(message[292]),
    .X(net214));
 sky130_fd_sc_hd__buf_1 input215 (.A(message[293]),
    .X(net215));
 sky130_fd_sc_hd__buf_1 input216 (.A(message[294]),
    .X(net216));
 sky130_fd_sc_hd__buf_1 input217 (.A(message[295]),
    .X(net217));
 sky130_fd_sc_hd__buf_1 input218 (.A(message[296]),
    .X(net218));
 sky130_fd_sc_hd__buf_1 input219 (.A(message[297]),
    .X(net219));
 sky130_fd_sc_hd__buf_1 input220 (.A(message[298]),
    .X(net220));
 sky130_fd_sc_hd__buf_1 input221 (.A(message[299]),
    .X(net221));
 sky130_fd_sc_hd__buf_1 input222 (.A(message[29]),
    .X(net222));
 sky130_fd_sc_hd__buf_1 input223 (.A(message[2]),
    .X(net223));
 sky130_fd_sc_hd__buf_1 input224 (.A(message[300]),
    .X(net224));
 sky130_fd_sc_hd__buf_1 input225 (.A(message[301]),
    .X(net225));
 sky130_fd_sc_hd__buf_1 input226 (.A(message[302]),
    .X(net226));
 sky130_fd_sc_hd__buf_1 input227 (.A(message[303]),
    .X(net227));
 sky130_fd_sc_hd__buf_1 input228 (.A(message[304]),
    .X(net228));
 sky130_fd_sc_hd__buf_1 input229 (.A(message[305]),
    .X(net229));
 sky130_fd_sc_hd__buf_1 input230 (.A(message[306]),
    .X(net230));
 sky130_fd_sc_hd__buf_1 input231 (.A(message[307]),
    .X(net231));
 sky130_fd_sc_hd__buf_1 input232 (.A(message[308]),
    .X(net232));
 sky130_fd_sc_hd__buf_1 input233 (.A(message[309]),
    .X(net233));
 sky130_fd_sc_hd__buf_1 input234 (.A(message[30]),
    .X(net234));
 sky130_fd_sc_hd__buf_1 input235 (.A(message[310]),
    .X(net235));
 sky130_fd_sc_hd__buf_1 input236 (.A(message[311]),
    .X(net236));
 sky130_fd_sc_hd__buf_1 input237 (.A(message[312]),
    .X(net237));
 sky130_fd_sc_hd__buf_1 input238 (.A(message[313]),
    .X(net238));
 sky130_fd_sc_hd__buf_1 input239 (.A(message[314]),
    .X(net239));
 sky130_fd_sc_hd__buf_1 input240 (.A(message[315]),
    .X(net240));
 sky130_fd_sc_hd__buf_1 input241 (.A(message[316]),
    .X(net241));
 sky130_fd_sc_hd__buf_1 input242 (.A(message[317]),
    .X(net242));
 sky130_fd_sc_hd__buf_1 input243 (.A(message[318]),
    .X(net243));
 sky130_fd_sc_hd__buf_1 input244 (.A(message[319]),
    .X(net244));
 sky130_fd_sc_hd__buf_1 input245 (.A(message[31]),
    .X(net245));
 sky130_fd_sc_hd__buf_1 input246 (.A(message[320]),
    .X(net246));
 sky130_fd_sc_hd__buf_1 input247 (.A(message[321]),
    .X(net247));
 sky130_fd_sc_hd__buf_1 input248 (.A(message[322]),
    .X(net248));
 sky130_fd_sc_hd__buf_1 input249 (.A(message[323]),
    .X(net249));
 sky130_fd_sc_hd__buf_1 input250 (.A(message[324]),
    .X(net250));
 sky130_fd_sc_hd__buf_1 input251 (.A(message[325]),
    .X(net251));
 sky130_fd_sc_hd__buf_1 input252 (.A(message[326]),
    .X(net252));
 sky130_fd_sc_hd__buf_1 input253 (.A(message[327]),
    .X(net253));
 sky130_fd_sc_hd__buf_1 input254 (.A(message[328]),
    .X(net254));
 sky130_fd_sc_hd__buf_1 input255 (.A(message[329]),
    .X(net255));
 sky130_fd_sc_hd__buf_1 input256 (.A(message[32]),
    .X(net256));
 sky130_fd_sc_hd__buf_1 input257 (.A(message[330]),
    .X(net257));
 sky130_fd_sc_hd__buf_1 input258 (.A(message[331]),
    .X(net258));
 sky130_fd_sc_hd__buf_1 input259 (.A(message[332]),
    .X(net259));
 sky130_fd_sc_hd__buf_1 input260 (.A(message[333]),
    .X(net260));
 sky130_fd_sc_hd__buf_1 input261 (.A(message[334]),
    .X(net261));
 sky130_fd_sc_hd__buf_1 input262 (.A(message[335]),
    .X(net262));
 sky130_fd_sc_hd__buf_1 input263 (.A(message[336]),
    .X(net263));
 sky130_fd_sc_hd__buf_1 input264 (.A(message[337]),
    .X(net264));
 sky130_fd_sc_hd__buf_1 input265 (.A(message[338]),
    .X(net265));
 sky130_fd_sc_hd__buf_1 input266 (.A(message[339]),
    .X(net266));
 sky130_fd_sc_hd__buf_1 input267 (.A(message[33]),
    .X(net267));
 sky130_fd_sc_hd__buf_1 input268 (.A(message[340]),
    .X(net268));
 sky130_fd_sc_hd__buf_1 input269 (.A(message[341]),
    .X(net269));
 sky130_fd_sc_hd__buf_1 input270 (.A(message[342]),
    .X(net270));
 sky130_fd_sc_hd__buf_1 input271 (.A(message[343]),
    .X(net271));
 sky130_fd_sc_hd__buf_1 input272 (.A(message[344]),
    .X(net272));
 sky130_fd_sc_hd__buf_1 input273 (.A(message[345]),
    .X(net273));
 sky130_fd_sc_hd__buf_1 input274 (.A(message[346]),
    .X(net274));
 sky130_fd_sc_hd__buf_1 input275 (.A(message[347]),
    .X(net275));
 sky130_fd_sc_hd__buf_1 input276 (.A(message[348]),
    .X(net276));
 sky130_fd_sc_hd__buf_1 input277 (.A(message[349]),
    .X(net277));
 sky130_fd_sc_hd__buf_1 input278 (.A(message[34]),
    .X(net278));
 sky130_fd_sc_hd__buf_1 input279 (.A(message[350]),
    .X(net279));
 sky130_fd_sc_hd__buf_1 input280 (.A(message[351]),
    .X(net280));
 sky130_fd_sc_hd__buf_1 input281 (.A(message[352]),
    .X(net281));
 sky130_fd_sc_hd__buf_1 input282 (.A(message[353]),
    .X(net282));
 sky130_fd_sc_hd__buf_1 input283 (.A(message[354]),
    .X(net283));
 sky130_fd_sc_hd__buf_1 input284 (.A(message[355]),
    .X(net284));
 sky130_fd_sc_hd__buf_1 input285 (.A(message[356]),
    .X(net552));
 sky130_fd_sc_hd__buf_1 input286 (.A(message[357]),
    .X(net553));
 sky130_fd_sc_hd__buf_1 input287 (.A(message[358]),
    .X(net554));
 sky130_fd_sc_hd__buf_1 input288 (.A(message[359]),
    .X(net555));
 sky130_fd_sc_hd__buf_1 input289 (.A(message[35]),
    .X(net556));
 sky130_fd_sc_hd__buf_1 input290 (.A(message[360]),
    .X(net557));
 sky130_fd_sc_hd__buf_1 input291 (.A(message[361]),
    .X(net558));
 sky130_fd_sc_hd__buf_1 input292 (.A(message[362]),
    .X(net559));
 sky130_fd_sc_hd__buf_1 input293 (.A(message[363]),
    .X(net560));
 sky130_fd_sc_hd__buf_1 input294 (.A(message[364]),
    .X(net561));
 sky130_fd_sc_hd__buf_1 input295 (.A(message[365]),
    .X(net562));
 sky130_fd_sc_hd__buf_1 input296 (.A(message[366]),
    .X(net563));
 sky130_fd_sc_hd__buf_1 input297 (.A(message[367]),
    .X(net564));
 sky130_fd_sc_hd__buf_1 input298 (.A(message[368]),
    .X(net565));
 sky130_fd_sc_hd__buf_1 input299 (.A(message[369]),
    .X(net566));
 sky130_fd_sc_hd__buf_1 input300 (.A(message[36]),
    .X(net567));
 sky130_fd_sc_hd__buf_1 input301 (.A(message[370]),
    .X(net568));
 sky130_fd_sc_hd__buf_1 input302 (.A(message[371]),
    .X(net569));
 sky130_fd_sc_hd__buf_1 input303 (.A(message[372]),
    .X(net570));
 sky130_fd_sc_hd__buf_1 input304 (.A(message[373]),
    .X(net571));
 sky130_fd_sc_hd__buf_1 input305 (.A(message[374]),
    .X(net572));
 sky130_fd_sc_hd__buf_1 input306 (.A(message[375]),
    .X(net573));
 sky130_fd_sc_hd__buf_1 input307 (.A(message[376]),
    .X(net574));
 sky130_fd_sc_hd__buf_1 input308 (.A(message[377]),
    .X(net575));
 sky130_fd_sc_hd__buf_1 input309 (.A(message[378]),
    .X(net576));
 sky130_fd_sc_hd__buf_1 input310 (.A(message[379]),
    .X(net577));
 sky130_fd_sc_hd__buf_1 input311 (.A(message[37]),
    .X(net578));
 sky130_fd_sc_hd__buf_1 input312 (.A(message[380]),
    .X(net579));
 sky130_fd_sc_hd__buf_1 input313 (.A(message[381]),
    .X(net580));
 sky130_fd_sc_hd__buf_1 input314 (.A(message[382]),
    .X(net581));
 sky130_fd_sc_hd__buf_1 input315 (.A(message[383]),
    .X(net582));
 sky130_fd_sc_hd__buf_1 input316 (.A(message[384]),
    .X(net583));
 sky130_fd_sc_hd__buf_1 input317 (.A(message[385]),
    .X(net584));
 sky130_fd_sc_hd__buf_1 input318 (.A(message[386]),
    .X(net585));
 sky130_fd_sc_hd__buf_1 input319 (.A(message[387]),
    .X(net586));
 sky130_fd_sc_hd__buf_1 input320 (.A(message[388]),
    .X(net587));
 sky130_fd_sc_hd__buf_1 input321 (.A(message[389]),
    .X(net588));
 sky130_fd_sc_hd__buf_1 input322 (.A(message[38]),
    .X(net589));
 sky130_fd_sc_hd__buf_1 input323 (.A(message[390]),
    .X(net590));
 sky130_fd_sc_hd__buf_1 input324 (.A(message[391]),
    .X(net591));
 sky130_fd_sc_hd__buf_1 input325 (.A(message[392]),
    .X(net592));
 sky130_fd_sc_hd__buf_1 input326 (.A(message[393]),
    .X(net593));
 sky130_fd_sc_hd__buf_1 input327 (.A(message[394]),
    .X(net594));
 sky130_fd_sc_hd__buf_1 input328 (.A(message[395]),
    .X(net595));
 sky130_fd_sc_hd__buf_1 input329 (.A(message[396]),
    .X(net596));
 sky130_fd_sc_hd__buf_1 input330 (.A(message[397]),
    .X(net597));
 sky130_fd_sc_hd__buf_1 input331 (.A(message[398]),
    .X(net598));
 sky130_fd_sc_hd__buf_1 input332 (.A(message[399]),
    .X(net599));
 sky130_fd_sc_hd__buf_1 input333 (.A(message[39]),
    .X(net600));
 sky130_fd_sc_hd__buf_1 input334 (.A(message[3]),
    .X(net601));
 sky130_fd_sc_hd__buf_1 input335 (.A(message[400]),
    .X(net602));
 sky130_fd_sc_hd__buf_1 input336 (.A(message[401]),
    .X(net603));
 sky130_fd_sc_hd__buf_1 input337 (.A(message[402]),
    .X(net604));
 sky130_fd_sc_hd__buf_1 input338 (.A(message[403]),
    .X(net605));
 sky130_fd_sc_hd__buf_1 input339 (.A(message[404]),
    .X(net606));
 sky130_fd_sc_hd__buf_1 input340 (.A(message[405]),
    .X(net607));
 sky130_fd_sc_hd__buf_1 input341 (.A(message[406]),
    .X(net608));
 sky130_fd_sc_hd__buf_1 input342 (.A(message[407]),
    .X(net609));
 sky130_fd_sc_hd__buf_1 input343 (.A(message[408]),
    .X(net610));
 sky130_fd_sc_hd__buf_1 input344 (.A(message[409]),
    .X(net611));
 sky130_fd_sc_hd__buf_1 input345 (.A(message[40]),
    .X(net612));
 sky130_fd_sc_hd__buf_1 input346 (.A(message[410]),
    .X(net613));
 sky130_fd_sc_hd__buf_1 input347 (.A(message[411]),
    .X(net614));
 sky130_fd_sc_hd__buf_1 input348 (.A(message[412]),
    .X(net615));
 sky130_fd_sc_hd__buf_1 input349 (.A(message[413]),
    .X(net616));
 sky130_fd_sc_hd__buf_1 input350 (.A(message[414]),
    .X(net617));
 sky130_fd_sc_hd__buf_1 input351 (.A(message[415]),
    .X(net618));
 sky130_fd_sc_hd__buf_1 input352 (.A(message[416]),
    .X(net619));
 sky130_fd_sc_hd__buf_1 input353 (.A(message[417]),
    .X(net620));
 sky130_fd_sc_hd__buf_1 input354 (.A(message[418]),
    .X(net621));
 sky130_fd_sc_hd__buf_1 input355 (.A(message[419]),
    .X(net622));
 sky130_fd_sc_hd__buf_1 input356 (.A(message[41]),
    .X(net623));
 sky130_fd_sc_hd__buf_1 input357 (.A(message[420]),
    .X(net624));
 sky130_fd_sc_hd__buf_1 input358 (.A(message[421]),
    .X(net625));
 sky130_fd_sc_hd__buf_1 input359 (.A(message[422]),
    .X(net626));
 sky130_fd_sc_hd__buf_1 input360 (.A(message[423]),
    .X(net627));
 sky130_fd_sc_hd__buf_1 input361 (.A(message[424]),
    .X(net628));
 sky130_fd_sc_hd__buf_1 input362 (.A(message[425]),
    .X(net629));
 sky130_fd_sc_hd__buf_1 input363 (.A(message[426]),
    .X(net630));
 sky130_fd_sc_hd__buf_1 input364 (.A(message[427]),
    .X(net631));
 sky130_fd_sc_hd__buf_1 input365 (.A(message[428]),
    .X(net632));
 sky130_fd_sc_hd__buf_1 input366 (.A(message[429]),
    .X(net633));
 sky130_fd_sc_hd__buf_1 input367 (.A(message[42]),
    .X(net634));
 sky130_fd_sc_hd__buf_1 input368 (.A(message[430]),
    .X(net635));
 sky130_fd_sc_hd__buf_1 input369 (.A(message[431]),
    .X(net636));
 sky130_fd_sc_hd__buf_1 input370 (.A(message[432]),
    .X(net637));
 sky130_fd_sc_hd__buf_1 input371 (.A(message[433]),
    .X(net638));
 sky130_fd_sc_hd__buf_1 input372 (.A(message[434]),
    .X(net639));
 sky130_fd_sc_hd__buf_1 input373 (.A(message[435]),
    .X(net640));
 sky130_fd_sc_hd__buf_1 input374 (.A(message[436]),
    .X(net641));
 sky130_fd_sc_hd__buf_1 input375 (.A(message[437]),
    .X(net642));
 sky130_fd_sc_hd__buf_1 input376 (.A(message[438]),
    .X(net643));
 sky130_fd_sc_hd__buf_1 input377 (.A(message[439]),
    .X(net644));
 sky130_fd_sc_hd__buf_1 input378 (.A(message[43]),
    .X(net645));
 sky130_fd_sc_hd__buf_1 input379 (.A(message[440]),
    .X(net646));
 sky130_fd_sc_hd__buf_1 input380 (.A(message[441]),
    .X(net647));
 sky130_fd_sc_hd__buf_1 input381 (.A(message[442]),
    .X(net648));
 sky130_fd_sc_hd__buf_1 input382 (.A(message[443]),
    .X(net649));
 sky130_fd_sc_hd__buf_1 input383 (.A(message[444]),
    .X(net650));
 sky130_fd_sc_hd__buf_1 input384 (.A(message[445]),
    .X(net651));
 sky130_fd_sc_hd__buf_1 input385 (.A(message[446]),
    .X(net652));
 sky130_fd_sc_hd__buf_1 input386 (.A(message[447]),
    .X(net653));
 sky130_fd_sc_hd__buf_1 input387 (.A(message[448]),
    .X(net654));
 sky130_fd_sc_hd__buf_1 input388 (.A(message[449]),
    .X(net655));
 sky130_fd_sc_hd__buf_1 input389 (.A(message[44]),
    .X(net656));
 sky130_fd_sc_hd__buf_1 input390 (.A(message[450]),
    .X(net657));
 sky130_fd_sc_hd__buf_1 input391 (.A(message[451]),
    .X(net658));
 sky130_fd_sc_hd__buf_1 input392 (.A(message[452]),
    .X(net659));
 sky130_fd_sc_hd__buf_1 input393 (.A(message[453]),
    .X(net660));
 sky130_fd_sc_hd__buf_1 input394 (.A(message[454]),
    .X(net661));
 sky130_fd_sc_hd__buf_1 input395 (.A(message[455]),
    .X(net662));
 sky130_fd_sc_hd__buf_1 input396 (.A(message[456]),
    .X(net663));
 sky130_fd_sc_hd__buf_1 input397 (.A(message[457]),
    .X(net664));
 sky130_fd_sc_hd__buf_1 input398 (.A(message[458]),
    .X(net665));
 sky130_fd_sc_hd__buf_1 input399 (.A(message[459]),
    .X(net666));
 sky130_fd_sc_hd__buf_1 input400 (.A(message[45]),
    .X(net667));
 sky130_fd_sc_hd__buf_1 input401 (.A(message[460]),
    .X(net668));
 sky130_fd_sc_hd__buf_1 input402 (.A(message[461]),
    .X(net669));
 sky130_fd_sc_hd__buf_1 input403 (.A(message[462]),
    .X(net670));
 sky130_fd_sc_hd__buf_1 input404 (.A(message[463]),
    .X(net671));
 sky130_fd_sc_hd__buf_1 input405 (.A(message[464]),
    .X(net672));
 sky130_fd_sc_hd__buf_1 input406 (.A(message[465]),
    .X(net673));
 sky130_fd_sc_hd__buf_1 input407 (.A(message[466]),
    .X(net674));
 sky130_fd_sc_hd__buf_1 input408 (.A(message[467]),
    .X(net675));
 sky130_fd_sc_hd__buf_1 input409 (.A(message[468]),
    .X(net676));
 sky130_fd_sc_hd__buf_1 input410 (.A(message[469]),
    .X(net677));
 sky130_fd_sc_hd__buf_1 input411 (.A(message[46]),
    .X(net678));
 sky130_fd_sc_hd__buf_1 input412 (.A(message[470]),
    .X(net679));
 sky130_fd_sc_hd__buf_1 input413 (.A(message[471]),
    .X(net680));
 sky130_fd_sc_hd__buf_1 input414 (.A(message[472]),
    .X(net681));
 sky130_fd_sc_hd__buf_1 input415 (.A(message[473]),
    .X(net682));
 sky130_fd_sc_hd__buf_1 input416 (.A(message[474]),
    .X(net683));
 sky130_fd_sc_hd__buf_1 input417 (.A(message[475]),
    .X(net684));
 sky130_fd_sc_hd__buf_1 input418 (.A(message[476]),
    .X(net685));
 sky130_fd_sc_hd__buf_1 input419 (.A(message[477]),
    .X(net686));
 sky130_fd_sc_hd__buf_1 input420 (.A(message[478]),
    .X(net687));
 sky130_fd_sc_hd__buf_1 input421 (.A(message[479]),
    .X(net688));
 sky130_fd_sc_hd__buf_1 input422 (.A(message[47]),
    .X(net689));
 sky130_fd_sc_hd__buf_1 input423 (.A(message[480]),
    .X(net690));
 sky130_fd_sc_hd__buf_1 input424 (.A(message[481]),
    .X(net691));
 sky130_fd_sc_hd__buf_1 input425 (.A(message[482]),
    .X(net692));
 sky130_fd_sc_hd__buf_1 input426 (.A(message[483]),
    .X(net693));
 sky130_fd_sc_hd__buf_1 input427 (.A(message[484]),
    .X(net694));
 sky130_fd_sc_hd__buf_1 input428 (.A(message[485]),
    .X(net695));
 sky130_fd_sc_hd__buf_1 input429 (.A(message[486]),
    .X(net696));
 sky130_fd_sc_hd__buf_1 input430 (.A(message[487]),
    .X(net697));
 sky130_fd_sc_hd__buf_1 input431 (.A(message[488]),
    .X(net698));
 sky130_fd_sc_hd__buf_1 input432 (.A(message[489]),
    .X(net699));
 sky130_fd_sc_hd__buf_1 input433 (.A(message[48]),
    .X(net700));
 sky130_fd_sc_hd__buf_1 input434 (.A(message[490]),
    .X(net701));
 sky130_fd_sc_hd__buf_1 input435 (.A(message[491]),
    .X(net702));
 sky130_fd_sc_hd__buf_1 input436 (.A(message[492]),
    .X(net703));
 sky130_fd_sc_hd__buf_1 input437 (.A(message[493]),
    .X(net704));
 sky130_fd_sc_hd__buf_1 input438 (.A(message[494]),
    .X(net705));
 sky130_fd_sc_hd__buf_1 input439 (.A(message[495]),
    .X(net706));
 sky130_fd_sc_hd__buf_1 input440 (.A(message[496]),
    .X(net707));
 sky130_fd_sc_hd__buf_1 input441 (.A(message[497]),
    .X(net708));
 sky130_fd_sc_hd__buf_1 input442 (.A(message[498]),
    .X(net709));
 sky130_fd_sc_hd__buf_1 input443 (.A(message[499]),
    .X(net710));
 sky130_fd_sc_hd__buf_1 input444 (.A(message[49]),
    .X(net711));
 sky130_fd_sc_hd__buf_1 input445 (.A(message[4]),
    .X(net712));
 sky130_fd_sc_hd__buf_1 input446 (.A(message[500]),
    .X(net713));
 sky130_fd_sc_hd__buf_1 input447 (.A(message[501]),
    .X(net714));
 sky130_fd_sc_hd__buf_1 input448 (.A(message[502]),
    .X(net715));
 sky130_fd_sc_hd__buf_1 input449 (.A(message[503]),
    .X(net716));
 sky130_fd_sc_hd__buf_1 input450 (.A(message[504]),
    .X(net717));
 sky130_fd_sc_hd__buf_1 input451 (.A(message[505]),
    .X(net718));
 sky130_fd_sc_hd__buf_1 input452 (.A(message[506]),
    .X(net719));
 sky130_fd_sc_hd__buf_1 input453 (.A(message[507]),
    .X(net720));
 sky130_fd_sc_hd__buf_1 input454 (.A(message[508]),
    .X(net721));
 sky130_fd_sc_hd__buf_1 input455 (.A(message[509]),
    .X(net722));
 sky130_fd_sc_hd__buf_1 input456 (.A(message[50]),
    .X(net723));
 sky130_fd_sc_hd__buf_1 input457 (.A(message[510]),
    .X(net724));
 sky130_fd_sc_hd__buf_1 input458 (.A(message[511]),
    .X(net725));
 sky130_fd_sc_hd__buf_1 input459 (.A(message[51]),
    .X(net726));
 sky130_fd_sc_hd__buf_1 input460 (.A(message[52]),
    .X(net727));
 sky130_fd_sc_hd__buf_1 input461 (.A(message[53]),
    .X(net728));
 sky130_fd_sc_hd__buf_1 input462 (.A(message[54]),
    .X(net729));
 sky130_fd_sc_hd__buf_1 input463 (.A(message[55]),
    .X(net730));
 sky130_fd_sc_hd__buf_1 input464 (.A(message[56]),
    .X(net731));
 sky130_fd_sc_hd__buf_1 input465 (.A(message[57]),
    .X(net732));
 sky130_fd_sc_hd__buf_1 input466 (.A(message[58]),
    .X(net733));
 sky130_fd_sc_hd__buf_1 input467 (.A(message[59]),
    .X(net734));
 sky130_fd_sc_hd__buf_1 input468 (.A(message[5]),
    .X(net735));
 sky130_fd_sc_hd__buf_1 input469 (.A(message[60]),
    .X(net736));
 sky130_fd_sc_hd__buf_1 input470 (.A(message[61]),
    .X(net737));
 sky130_fd_sc_hd__buf_1 input471 (.A(message[62]),
    .X(net738));
 sky130_fd_sc_hd__buf_1 input472 (.A(message[63]),
    .X(net739));
 sky130_fd_sc_hd__buf_1 input473 (.A(message[64]),
    .X(net740));
 sky130_fd_sc_hd__buf_1 input474 (.A(message[65]),
    .X(net741));
 sky130_fd_sc_hd__buf_1 input475 (.A(message[66]),
    .X(net742));
 sky130_fd_sc_hd__buf_1 input476 (.A(message[67]),
    .X(net743));
 sky130_fd_sc_hd__buf_1 input477 (.A(message[68]),
    .X(net744));
 sky130_fd_sc_hd__buf_1 input478 (.A(message[69]),
    .X(net745));
 sky130_fd_sc_hd__buf_1 input479 (.A(message[6]),
    .X(net746));
 sky130_fd_sc_hd__buf_1 input480 (.A(message[70]),
    .X(net747));
 sky130_fd_sc_hd__buf_1 input481 (.A(message[71]),
    .X(net748));
 sky130_fd_sc_hd__buf_1 input482 (.A(message[72]),
    .X(net749));
 sky130_fd_sc_hd__buf_1 input483 (.A(message[73]),
    .X(net750));
 sky130_fd_sc_hd__buf_1 input484 (.A(message[74]),
    .X(net751));
 sky130_fd_sc_hd__buf_1 input485 (.A(message[75]),
    .X(net752));
 sky130_fd_sc_hd__buf_1 input486 (.A(message[76]),
    .X(net753));
 sky130_fd_sc_hd__buf_1 input487 (.A(message[77]),
    .X(net754));
 sky130_fd_sc_hd__buf_1 input488 (.A(message[78]),
    .X(net755));
 sky130_fd_sc_hd__buf_1 input489 (.A(message[79]),
    .X(net756));
 sky130_fd_sc_hd__buf_1 input490 (.A(message[7]),
    .X(net757));
 sky130_fd_sc_hd__buf_1 input491 (.A(message[80]),
    .X(net758));
 sky130_fd_sc_hd__buf_1 input492 (.A(message[81]),
    .X(net759));
 sky130_fd_sc_hd__buf_1 input493 (.A(message[82]),
    .X(net760));
 sky130_fd_sc_hd__buf_1 input494 (.A(message[83]),
    .X(net761));
 sky130_fd_sc_hd__buf_1 input495 (.A(message[84]),
    .X(net762));
 sky130_fd_sc_hd__buf_1 input496 (.A(message[85]),
    .X(net763));
 sky130_fd_sc_hd__buf_1 input497 (.A(message[86]),
    .X(net764));
 sky130_fd_sc_hd__buf_1 input498 (.A(message[87]),
    .X(net765));
 sky130_fd_sc_hd__buf_1 input499 (.A(message[88]),
    .X(net766));
 sky130_fd_sc_hd__buf_1 input500 (.A(message[89]),
    .X(net767));
 sky130_fd_sc_hd__buf_1 input501 (.A(message[8]),
    .X(net768));
 sky130_fd_sc_hd__buf_1 input502 (.A(message[90]),
    .X(net769));
 sky130_fd_sc_hd__buf_1 input503 (.A(message[91]),
    .X(net770));
 sky130_fd_sc_hd__buf_1 input504 (.A(message[92]),
    .X(net771));
 sky130_fd_sc_hd__buf_1 input505 (.A(message[93]),
    .X(net772));
 sky130_fd_sc_hd__buf_1 input506 (.A(message[94]),
    .X(net773));
 sky130_fd_sc_hd__buf_1 input507 (.A(message[95]),
    .X(net774));
 sky130_fd_sc_hd__buf_1 input508 (.A(message[96]),
    .X(net775));
 sky130_fd_sc_hd__buf_1 input509 (.A(message[97]),
    .X(net776));
 sky130_fd_sc_hd__buf_1 input510 (.A(message[98]),
    .X(net777));
 sky130_fd_sc_hd__buf_1 input511 (.A(message[99]),
    .X(net778));
 sky130_fd_sc_hd__buf_1 input512 (.A(message[9]),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_1 input513 (.A(reset),
    .X(net780));
 sky130_fd_sc_hd__buf_1 output514 (.A(net781),
    .X(hashvalue[0]));
 sky130_fd_sc_hd__buf_1 output515 (.A(net782),
    .X(hashvalue[100]));
 sky130_fd_sc_hd__buf_1 output516 (.A(net783),
    .X(hashvalue[101]));
 sky130_fd_sc_hd__buf_1 output517 (.A(net784),
    .X(hashvalue[102]));
 sky130_fd_sc_hd__buf_1 output518 (.A(net785),
    .X(hashvalue[103]));
 sky130_fd_sc_hd__buf_1 output519 (.A(net786),
    .X(hashvalue[104]));
 sky130_fd_sc_hd__buf_1 output520 (.A(net787),
    .X(hashvalue[105]));
 sky130_fd_sc_hd__buf_1 output521 (.A(net788),
    .X(hashvalue[106]));
 sky130_fd_sc_hd__buf_1 output522 (.A(net789),
    .X(hashvalue[107]));
 sky130_fd_sc_hd__buf_1 output523 (.A(net790),
    .X(hashvalue[108]));
 sky130_fd_sc_hd__buf_1 output524 (.A(net791),
    .X(hashvalue[109]));
 sky130_fd_sc_hd__buf_1 output525 (.A(net792),
    .X(hashvalue[10]));
 sky130_fd_sc_hd__buf_1 output526 (.A(net793),
    .X(hashvalue[110]));
 sky130_fd_sc_hd__buf_1 output527 (.A(net794),
    .X(hashvalue[111]));
 sky130_fd_sc_hd__buf_1 output528 (.A(net795),
    .X(hashvalue[112]));
 sky130_fd_sc_hd__buf_1 output529 (.A(net796),
    .X(hashvalue[113]));
 sky130_fd_sc_hd__buf_1 output530 (.A(net797),
    .X(hashvalue[114]));
 sky130_fd_sc_hd__buf_1 output531 (.A(net798),
    .X(hashvalue[115]));
 sky130_fd_sc_hd__buf_1 output532 (.A(net799),
    .X(hashvalue[116]));
 sky130_fd_sc_hd__buf_1 output533 (.A(net800),
    .X(hashvalue[117]));
 sky130_fd_sc_hd__buf_1 output534 (.A(net801),
    .X(hashvalue[118]));
 sky130_fd_sc_hd__buf_1 output535 (.A(net802),
    .X(hashvalue[119]));
 sky130_fd_sc_hd__buf_1 output536 (.A(net803),
    .X(hashvalue[11]));
 sky130_fd_sc_hd__buf_1 output537 (.A(net804),
    .X(hashvalue[120]));
 sky130_fd_sc_hd__buf_1 output538 (.A(net805),
    .X(hashvalue[121]));
 sky130_fd_sc_hd__buf_1 output539 (.A(net806),
    .X(hashvalue[122]));
 sky130_fd_sc_hd__buf_1 output540 (.A(net807),
    .X(hashvalue[123]));
 sky130_fd_sc_hd__buf_1 output541 (.A(net808),
    .X(hashvalue[124]));
 sky130_fd_sc_hd__buf_1 output542 (.A(net809),
    .X(hashvalue[125]));
 sky130_fd_sc_hd__buf_1 output543 (.A(net810),
    .X(hashvalue[126]));
 sky130_fd_sc_hd__buf_1 output544 (.A(net811),
    .X(hashvalue[127]));
 sky130_fd_sc_hd__buf_1 output545 (.A(net812),
    .X(hashvalue[128]));
 sky130_fd_sc_hd__buf_1 output546 (.A(net813),
    .X(hashvalue[129]));
 sky130_fd_sc_hd__buf_1 output547 (.A(net814),
    .X(hashvalue[12]));
 sky130_fd_sc_hd__buf_1 output548 (.A(net815),
    .X(hashvalue[130]));
 sky130_fd_sc_hd__buf_1 output549 (.A(net816),
    .X(hashvalue[131]));
 sky130_fd_sc_hd__buf_1 output550 (.A(net817),
    .X(hashvalue[132]));
 sky130_fd_sc_hd__buf_1 output551 (.A(net818),
    .X(hashvalue[133]));
 sky130_fd_sc_hd__buf_1 output552 (.A(net819),
    .X(hashvalue[134]));
 sky130_fd_sc_hd__buf_1 output553 (.A(net820),
    .X(hashvalue[135]));
 sky130_fd_sc_hd__buf_1 output554 (.A(net821),
    .X(hashvalue[136]));
 sky130_fd_sc_hd__buf_1 output555 (.A(net822),
    .X(hashvalue[137]));
 sky130_fd_sc_hd__buf_1 output556 (.A(net823),
    .X(hashvalue[138]));
 sky130_fd_sc_hd__buf_1 output557 (.A(net824),
    .X(hashvalue[139]));
 sky130_fd_sc_hd__buf_1 output558 (.A(net825),
    .X(hashvalue[13]));
 sky130_fd_sc_hd__buf_1 output559 (.A(net826),
    .X(hashvalue[140]));
 sky130_fd_sc_hd__buf_1 output560 (.A(net827),
    .X(hashvalue[141]));
 sky130_fd_sc_hd__buf_1 output561 (.A(net828),
    .X(hashvalue[142]));
 sky130_fd_sc_hd__buf_1 output562 (.A(net829),
    .X(hashvalue[143]));
 sky130_fd_sc_hd__buf_1 output563 (.A(net830),
    .X(hashvalue[144]));
 sky130_fd_sc_hd__buf_1 output564 (.A(net831),
    .X(hashvalue[145]));
 sky130_fd_sc_hd__buf_1 output565 (.A(net832),
    .X(hashvalue[146]));
 sky130_fd_sc_hd__buf_1 output566 (.A(net833),
    .X(hashvalue[147]));
 sky130_fd_sc_hd__buf_1 output567 (.A(net834),
    .X(hashvalue[148]));
 sky130_fd_sc_hd__buf_1 output568 (.A(net835),
    .X(hashvalue[149]));
 sky130_fd_sc_hd__buf_1 output569 (.A(net836),
    .X(hashvalue[14]));
 sky130_fd_sc_hd__buf_1 output570 (.A(net837),
    .X(hashvalue[150]));
 sky130_fd_sc_hd__buf_1 output571 (.A(net838),
    .X(hashvalue[151]));
 sky130_fd_sc_hd__buf_1 output572 (.A(net839),
    .X(hashvalue[152]));
 sky130_fd_sc_hd__buf_1 output573 (.A(net840),
    .X(hashvalue[153]));
 sky130_fd_sc_hd__buf_1 output574 (.A(net841),
    .X(hashvalue[154]));
 sky130_fd_sc_hd__buf_1 output575 (.A(net842),
    .X(hashvalue[155]));
 sky130_fd_sc_hd__buf_1 output576 (.A(net843),
    .X(hashvalue[156]));
 sky130_fd_sc_hd__buf_1 output577 (.A(net844),
    .X(hashvalue[157]));
 sky130_fd_sc_hd__buf_1 output578 (.A(net845),
    .X(hashvalue[158]));
 sky130_fd_sc_hd__buf_1 output579 (.A(net846),
    .X(hashvalue[159]));
 sky130_fd_sc_hd__buf_1 output580 (.A(net847),
    .X(hashvalue[15]));
 sky130_fd_sc_hd__buf_1 output581 (.A(net848),
    .X(hashvalue[160]));
 sky130_fd_sc_hd__buf_1 output582 (.A(net849),
    .X(hashvalue[161]));
 sky130_fd_sc_hd__buf_1 output583 (.A(net850),
    .X(hashvalue[162]));
 sky130_fd_sc_hd__buf_1 output584 (.A(net851),
    .X(hashvalue[163]));
 sky130_fd_sc_hd__buf_1 output585 (.A(net852),
    .X(hashvalue[164]));
 sky130_fd_sc_hd__buf_1 output586 (.A(net853),
    .X(hashvalue[165]));
 sky130_fd_sc_hd__buf_1 output587 (.A(net854),
    .X(hashvalue[166]));
 sky130_fd_sc_hd__buf_1 output588 (.A(net855),
    .X(hashvalue[167]));
 sky130_fd_sc_hd__buf_1 output589 (.A(net856),
    .X(hashvalue[168]));
 sky130_fd_sc_hd__buf_1 output590 (.A(net857),
    .X(hashvalue[169]));
 sky130_fd_sc_hd__buf_1 output591 (.A(net858),
    .X(hashvalue[16]));
 sky130_fd_sc_hd__buf_1 output592 (.A(net859),
    .X(hashvalue[170]));
 sky130_fd_sc_hd__buf_1 output593 (.A(net860),
    .X(hashvalue[171]));
 sky130_fd_sc_hd__buf_1 output594 (.A(net861),
    .X(hashvalue[172]));
 sky130_fd_sc_hd__buf_1 output595 (.A(net862),
    .X(hashvalue[173]));
 sky130_fd_sc_hd__buf_1 output596 (.A(net863),
    .X(hashvalue[174]));
 sky130_fd_sc_hd__buf_1 output597 (.A(net864),
    .X(hashvalue[175]));
 sky130_fd_sc_hd__buf_1 output598 (.A(net865),
    .X(hashvalue[176]));
 sky130_fd_sc_hd__buf_1 output599 (.A(net866),
    .X(hashvalue[177]));
 sky130_fd_sc_hd__buf_1 output600 (.A(net867),
    .X(hashvalue[178]));
 sky130_fd_sc_hd__buf_1 output601 (.A(net868),
    .X(hashvalue[179]));
 sky130_fd_sc_hd__buf_1 output602 (.A(net869),
    .X(hashvalue[17]));
 sky130_fd_sc_hd__buf_1 output603 (.A(net870),
    .X(hashvalue[180]));
 sky130_fd_sc_hd__buf_1 output604 (.A(net871),
    .X(hashvalue[181]));
 sky130_fd_sc_hd__buf_1 output605 (.A(net872),
    .X(hashvalue[182]));
 sky130_fd_sc_hd__buf_1 output606 (.A(net873),
    .X(hashvalue[183]));
 sky130_fd_sc_hd__buf_1 output607 (.A(net874),
    .X(hashvalue[184]));
 sky130_fd_sc_hd__buf_1 output608 (.A(net875),
    .X(hashvalue[185]));
 sky130_fd_sc_hd__buf_1 output609 (.A(net876),
    .X(hashvalue[186]));
 sky130_fd_sc_hd__buf_1 output610 (.A(net877),
    .X(hashvalue[187]));
 sky130_fd_sc_hd__buf_1 output611 (.A(net878),
    .X(hashvalue[188]));
 sky130_fd_sc_hd__buf_1 output612 (.A(net879),
    .X(hashvalue[189]));
 sky130_fd_sc_hd__buf_1 output613 (.A(net880),
    .X(hashvalue[18]));
 sky130_fd_sc_hd__buf_1 output614 (.A(net881),
    .X(hashvalue[190]));
 sky130_fd_sc_hd__buf_1 output615 (.A(net882),
    .X(hashvalue[191]));
 sky130_fd_sc_hd__buf_1 output616 (.A(net883),
    .X(hashvalue[192]));
 sky130_fd_sc_hd__buf_1 output617 (.A(net884),
    .X(hashvalue[193]));
 sky130_fd_sc_hd__buf_1 output618 (.A(net885),
    .X(hashvalue[194]));
 sky130_fd_sc_hd__buf_1 output619 (.A(net886),
    .X(hashvalue[195]));
 sky130_fd_sc_hd__buf_1 output620 (.A(net887),
    .X(hashvalue[196]));
 sky130_fd_sc_hd__buf_1 output621 (.A(net888),
    .X(hashvalue[197]));
 sky130_fd_sc_hd__buf_1 output622 (.A(net889),
    .X(hashvalue[198]));
 sky130_fd_sc_hd__buf_1 output623 (.A(net890),
    .X(hashvalue[199]));
 sky130_fd_sc_hd__buf_1 output624 (.A(net891),
    .X(hashvalue[19]));
 sky130_fd_sc_hd__buf_1 output625 (.A(net892),
    .X(hashvalue[1]));
 sky130_fd_sc_hd__buf_1 output626 (.A(net893),
    .X(hashvalue[200]));
 sky130_fd_sc_hd__buf_1 output627 (.A(net894),
    .X(hashvalue[201]));
 sky130_fd_sc_hd__buf_1 output628 (.A(net895),
    .X(hashvalue[202]));
 sky130_fd_sc_hd__buf_1 output629 (.A(net896),
    .X(hashvalue[203]));
 sky130_fd_sc_hd__buf_1 output630 (.A(net897),
    .X(hashvalue[204]));
 sky130_fd_sc_hd__buf_1 output631 (.A(net898),
    .X(hashvalue[205]));
 sky130_fd_sc_hd__buf_1 output632 (.A(net899),
    .X(hashvalue[206]));
 sky130_fd_sc_hd__buf_1 output633 (.A(net900),
    .X(hashvalue[207]));
 sky130_fd_sc_hd__buf_1 output634 (.A(net901),
    .X(hashvalue[208]));
 sky130_fd_sc_hd__buf_1 output635 (.A(net902),
    .X(hashvalue[209]));
 sky130_fd_sc_hd__buf_1 output636 (.A(net903),
    .X(hashvalue[20]));
 sky130_fd_sc_hd__buf_1 output637 (.A(net904),
    .X(hashvalue[210]));
 sky130_fd_sc_hd__buf_1 output638 (.A(net905),
    .X(hashvalue[211]));
 sky130_fd_sc_hd__buf_1 output639 (.A(net906),
    .X(hashvalue[212]));
 sky130_fd_sc_hd__buf_1 output640 (.A(net907),
    .X(hashvalue[213]));
 sky130_fd_sc_hd__buf_1 output641 (.A(net908),
    .X(hashvalue[214]));
 sky130_fd_sc_hd__buf_1 output642 (.A(net909),
    .X(hashvalue[215]));
 sky130_fd_sc_hd__buf_1 output643 (.A(net910),
    .X(hashvalue[216]));
 sky130_fd_sc_hd__buf_1 output644 (.A(net911),
    .X(hashvalue[217]));
 sky130_fd_sc_hd__buf_1 output645 (.A(net912),
    .X(hashvalue[218]));
 sky130_fd_sc_hd__buf_1 output646 (.A(net913),
    .X(hashvalue[219]));
 sky130_fd_sc_hd__buf_1 output647 (.A(net914),
    .X(hashvalue[21]));
 sky130_fd_sc_hd__buf_1 output648 (.A(net915),
    .X(hashvalue[220]));
 sky130_fd_sc_hd__buf_1 output649 (.A(net916),
    .X(hashvalue[221]));
 sky130_fd_sc_hd__buf_1 output650 (.A(net917),
    .X(hashvalue[222]));
 sky130_fd_sc_hd__buf_1 output651 (.A(net918),
    .X(hashvalue[223]));
 sky130_fd_sc_hd__buf_1 output652 (.A(net919),
    .X(hashvalue[224]));
 sky130_fd_sc_hd__buf_1 output653 (.A(net920),
    .X(hashvalue[225]));
 sky130_fd_sc_hd__buf_1 output654 (.A(net921),
    .X(hashvalue[226]));
 sky130_fd_sc_hd__buf_1 output655 (.A(net922),
    .X(hashvalue[227]));
 sky130_fd_sc_hd__buf_1 output656 (.A(net923),
    .X(hashvalue[228]));
 sky130_fd_sc_hd__buf_1 output657 (.A(net924),
    .X(hashvalue[229]));
 sky130_fd_sc_hd__buf_1 output658 (.A(net925),
    .X(hashvalue[22]));
 sky130_fd_sc_hd__buf_1 output659 (.A(net926),
    .X(hashvalue[230]));
 sky130_fd_sc_hd__buf_1 output660 (.A(net927),
    .X(hashvalue[231]));
 sky130_fd_sc_hd__buf_1 output661 (.A(net928),
    .X(hashvalue[232]));
 sky130_fd_sc_hd__buf_1 output662 (.A(net929),
    .X(hashvalue[233]));
 sky130_fd_sc_hd__buf_1 output663 (.A(net930),
    .X(hashvalue[234]));
 sky130_fd_sc_hd__buf_1 output664 (.A(net931),
    .X(hashvalue[235]));
 sky130_fd_sc_hd__buf_1 output665 (.A(net932),
    .X(hashvalue[236]));
 sky130_fd_sc_hd__buf_1 output666 (.A(net933),
    .X(hashvalue[237]));
 sky130_fd_sc_hd__buf_1 output667 (.A(net934),
    .X(hashvalue[238]));
 sky130_fd_sc_hd__buf_1 output668 (.A(net935),
    .X(hashvalue[239]));
 sky130_fd_sc_hd__buf_1 output669 (.A(net936),
    .X(hashvalue[23]));
 sky130_fd_sc_hd__buf_1 output670 (.A(net937),
    .X(hashvalue[240]));
 sky130_fd_sc_hd__buf_1 output671 (.A(net938),
    .X(hashvalue[241]));
 sky130_fd_sc_hd__buf_1 output672 (.A(net939),
    .X(hashvalue[242]));
 sky130_fd_sc_hd__buf_1 output673 (.A(net940),
    .X(hashvalue[243]));
 sky130_fd_sc_hd__buf_1 output674 (.A(net941),
    .X(hashvalue[244]));
 sky130_fd_sc_hd__buf_1 output675 (.A(net942),
    .X(hashvalue[245]));
 sky130_fd_sc_hd__buf_1 output676 (.A(net943),
    .X(hashvalue[246]));
 sky130_fd_sc_hd__buf_1 output677 (.A(net944),
    .X(hashvalue[247]));
 sky130_fd_sc_hd__buf_1 output678 (.A(net945),
    .X(hashvalue[248]));
 sky130_fd_sc_hd__buf_1 output679 (.A(net946),
    .X(hashvalue[249]));
 sky130_fd_sc_hd__buf_1 output680 (.A(net947),
    .X(hashvalue[24]));
 sky130_fd_sc_hd__buf_1 output681 (.A(net948),
    .X(hashvalue[250]));
 sky130_fd_sc_hd__buf_1 output682 (.A(net949),
    .X(hashvalue[251]));
 sky130_fd_sc_hd__buf_1 output683 (.A(net950),
    .X(hashvalue[252]));
 sky130_fd_sc_hd__buf_1 output684 (.A(net951),
    .X(hashvalue[253]));
 sky130_fd_sc_hd__buf_1 output685 (.A(net952),
    .X(hashvalue[254]));
 sky130_fd_sc_hd__buf_1 output686 (.A(net953),
    .X(hashvalue[255]));
 sky130_fd_sc_hd__buf_1 output687 (.A(net954),
    .X(hashvalue[25]));
 sky130_fd_sc_hd__buf_1 output688 (.A(net955),
    .X(hashvalue[26]));
 sky130_fd_sc_hd__buf_1 output689 (.A(net956),
    .X(hashvalue[27]));
 sky130_fd_sc_hd__buf_1 output690 (.A(net957),
    .X(hashvalue[28]));
 sky130_fd_sc_hd__buf_1 output691 (.A(net958),
    .X(hashvalue[29]));
 sky130_fd_sc_hd__buf_1 output692 (.A(net959),
    .X(hashvalue[2]));
 sky130_fd_sc_hd__buf_1 output693 (.A(net960),
    .X(hashvalue[30]));
 sky130_fd_sc_hd__buf_1 output694 (.A(net961),
    .X(hashvalue[31]));
 sky130_fd_sc_hd__buf_1 output695 (.A(net962),
    .X(hashvalue[32]));
 sky130_fd_sc_hd__buf_1 output696 (.A(net963),
    .X(hashvalue[33]));
 sky130_fd_sc_hd__buf_1 output697 (.A(net964),
    .X(hashvalue[34]));
 sky130_fd_sc_hd__buf_1 output698 (.A(net965),
    .X(hashvalue[35]));
 sky130_fd_sc_hd__buf_1 output699 (.A(net966),
    .X(hashvalue[36]));
 sky130_fd_sc_hd__buf_1 output700 (.A(net967),
    .X(hashvalue[37]));
 sky130_fd_sc_hd__buf_1 output701 (.A(net968),
    .X(hashvalue[38]));
 sky130_fd_sc_hd__buf_1 output702 (.A(net969),
    .X(hashvalue[39]));
 sky130_fd_sc_hd__buf_1 output703 (.A(net970),
    .X(hashvalue[3]));
 sky130_fd_sc_hd__buf_1 output704 (.A(net971),
    .X(hashvalue[40]));
 sky130_fd_sc_hd__buf_1 output705 (.A(net972),
    .X(hashvalue[41]));
 sky130_fd_sc_hd__buf_1 output706 (.A(net973),
    .X(hashvalue[42]));
 sky130_fd_sc_hd__buf_1 output707 (.A(net974),
    .X(hashvalue[43]));
 sky130_fd_sc_hd__buf_1 output708 (.A(net975),
    .X(hashvalue[44]));
 sky130_fd_sc_hd__buf_1 output709 (.A(net976),
    .X(hashvalue[45]));
 sky130_fd_sc_hd__buf_1 output710 (.A(net977),
    .X(hashvalue[46]));
 sky130_fd_sc_hd__buf_1 output711 (.A(net978),
    .X(hashvalue[47]));
 sky130_fd_sc_hd__buf_1 output712 (.A(net979),
    .X(hashvalue[48]));
 sky130_fd_sc_hd__buf_1 output713 (.A(net980),
    .X(hashvalue[49]));
 sky130_fd_sc_hd__buf_1 output714 (.A(net981),
    .X(hashvalue[4]));
 sky130_fd_sc_hd__buf_1 output715 (.A(net982),
    .X(hashvalue[50]));
 sky130_fd_sc_hd__buf_1 output716 (.A(net983),
    .X(hashvalue[51]));
 sky130_fd_sc_hd__buf_1 output717 (.A(net984),
    .X(hashvalue[52]));
 sky130_fd_sc_hd__buf_1 output718 (.A(net985),
    .X(hashvalue[53]));
 sky130_fd_sc_hd__buf_1 output719 (.A(net986),
    .X(hashvalue[54]));
 sky130_fd_sc_hd__buf_1 output720 (.A(net987),
    .X(hashvalue[55]));
 sky130_fd_sc_hd__buf_1 output721 (.A(net988),
    .X(hashvalue[56]));
 sky130_fd_sc_hd__buf_1 output722 (.A(net989),
    .X(hashvalue[57]));
 sky130_fd_sc_hd__buf_1 output723 (.A(net990),
    .X(hashvalue[58]));
 sky130_fd_sc_hd__buf_1 output724 (.A(net991),
    .X(hashvalue[59]));
 sky130_fd_sc_hd__buf_1 output725 (.A(net992),
    .X(hashvalue[5]));
 sky130_fd_sc_hd__buf_1 output726 (.A(net993),
    .X(hashvalue[60]));
 sky130_fd_sc_hd__buf_1 output727 (.A(net994),
    .X(hashvalue[61]));
 sky130_fd_sc_hd__buf_1 output728 (.A(net995),
    .X(hashvalue[62]));
 sky130_fd_sc_hd__buf_1 output729 (.A(net996),
    .X(hashvalue[63]));
 sky130_fd_sc_hd__buf_1 output730 (.A(net997),
    .X(hashvalue[64]));
 sky130_fd_sc_hd__buf_1 output731 (.A(net998),
    .X(hashvalue[65]));
 sky130_fd_sc_hd__buf_1 output732 (.A(net999),
    .X(hashvalue[66]));
 sky130_fd_sc_hd__buf_1 output733 (.A(net1000),
    .X(hashvalue[67]));
 sky130_fd_sc_hd__buf_1 output734 (.A(net1001),
    .X(hashvalue[68]));
 sky130_fd_sc_hd__buf_1 output735 (.A(net1002),
    .X(hashvalue[69]));
 sky130_fd_sc_hd__buf_1 output736 (.A(net1003),
    .X(hashvalue[6]));
 sky130_fd_sc_hd__buf_1 output737 (.A(net1004),
    .X(hashvalue[70]));
 sky130_fd_sc_hd__buf_1 output738 (.A(net1005),
    .X(hashvalue[71]));
 sky130_fd_sc_hd__buf_1 output739 (.A(net1006),
    .X(hashvalue[72]));
 sky130_fd_sc_hd__buf_1 output740 (.A(net1007),
    .X(hashvalue[73]));
 sky130_fd_sc_hd__buf_1 output741 (.A(net1008),
    .X(hashvalue[74]));
 sky130_fd_sc_hd__buf_1 output742 (.A(net1009),
    .X(hashvalue[75]));
 sky130_fd_sc_hd__buf_1 output743 (.A(net1010),
    .X(hashvalue[76]));
 sky130_fd_sc_hd__buf_1 output744 (.A(net1011),
    .X(hashvalue[77]));
 sky130_fd_sc_hd__buf_1 output745 (.A(net1012),
    .X(hashvalue[78]));
 sky130_fd_sc_hd__buf_1 output746 (.A(net1013),
    .X(hashvalue[79]));
 sky130_fd_sc_hd__buf_1 output747 (.A(net1014),
    .X(hashvalue[7]));
 sky130_fd_sc_hd__buf_1 output748 (.A(net1015),
    .X(hashvalue[80]));
 sky130_fd_sc_hd__buf_1 output749 (.A(net1016),
    .X(hashvalue[81]));
 sky130_fd_sc_hd__buf_1 output750 (.A(net1017),
    .X(hashvalue[82]));
 sky130_fd_sc_hd__buf_1 output751 (.A(net1018),
    .X(hashvalue[83]));
 sky130_fd_sc_hd__buf_1 output752 (.A(net1019),
    .X(hashvalue[84]));
 sky130_fd_sc_hd__buf_1 output753 (.A(net1020),
    .X(hashvalue[85]));
 sky130_fd_sc_hd__buf_1 output754 (.A(net1021),
    .X(hashvalue[86]));
 sky130_fd_sc_hd__buf_1 output755 (.A(net1022),
    .X(hashvalue[87]));
 sky130_fd_sc_hd__buf_1 output756 (.A(net1023),
    .X(hashvalue[88]));
 sky130_fd_sc_hd__buf_1 output757 (.A(net1024),
    .X(hashvalue[89]));
 sky130_fd_sc_hd__buf_1 output758 (.A(net1025),
    .X(hashvalue[8]));
 sky130_fd_sc_hd__buf_1 output759 (.A(net1026),
    .X(hashvalue[90]));
 sky130_fd_sc_hd__buf_1 output760 (.A(net1027),
    .X(hashvalue[91]));
 sky130_fd_sc_hd__buf_1 output761 (.A(net1028),
    .X(hashvalue[92]));
 sky130_fd_sc_hd__buf_1 output762 (.A(net1029),
    .X(hashvalue[93]));
 sky130_fd_sc_hd__buf_1 output763 (.A(net1030),
    .X(hashvalue[94]));
 sky130_fd_sc_hd__buf_1 output764 (.A(net1031),
    .X(hashvalue[95]));
 sky130_fd_sc_hd__buf_1 output765 (.A(net1032),
    .X(hashvalue[96]));
 sky130_fd_sc_hd__buf_1 output766 (.A(net1033),
    .X(hashvalue[97]));
 sky130_fd_sc_hd__buf_1 output767 (.A(net1034),
    .X(hashvalue[98]));
 sky130_fd_sc_hd__buf_1 output768 (.A(net1035),
    .X(hashvalue[99]));
 sky130_fd_sc_hd__buf_1 output769 (.A(net1036),
    .X(hashvalue[9]));
 sky130_fd_sc_hd__buf_1 output770 (.A(net1037),
    .X(ready));
 sky130_fd_sc_hd__clkbuf_1 load_slew771 (.A(net1039),
    .X(net1038));
 sky130_fd_sc_hd__clkbuf_1 load_slew772 (.A(net780),
    .X(net1039));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_147_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_193_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_194_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_198_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_199_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_200_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_201_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_202_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_203_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_204_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_205_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_206_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_207_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_208_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_209_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_210_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_211_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_212_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_213_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_214_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_215_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_216_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_217_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_218_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_218_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_219_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_219_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_220_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_220_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_221_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_222_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_223_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_224_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_225_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_226_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_227_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_227_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_228_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_229_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_230_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_230_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_231_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_232_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_232_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_233_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_234_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_234_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_235_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_235_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_236_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_236_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_237_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_238_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_239_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_240_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_241_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_242_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_243_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_244_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_244_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_245_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_245_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_246_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_246_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_247_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_247_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_248_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_248_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_249_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_249_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_250_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_250_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_251_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_251_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_252_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_252_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_253_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_253_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_254_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_254_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_255_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_255_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_256_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_256_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_257_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_257_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_258_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_258_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_259_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_259_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_260_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_260_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_261_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_261_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_262_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_262_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_263_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_263_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_264_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_264_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_265_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_265_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_266_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_266_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_267_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_267_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_268_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_268_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_269_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_269_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_270_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_270_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_271_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_271_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_272_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_272_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_273_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_273_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_274_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_274_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_275_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_275_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_276_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_276_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_277_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_277_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_278_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_278_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_279_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_279_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_280_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_280_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_281_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_281_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_282_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_282_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_283_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_283_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_284_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_284_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_285_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_285_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_286_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_286_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_287_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_287_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_288_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_288_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_289_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_289_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_290_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_290_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_0__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_1__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_2__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_3__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_4__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_5__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_6__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_7__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_5_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_8__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_8__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_9__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_9__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_10__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_10__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_11__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_11__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_12__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_12__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_13__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_13__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_14__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_14__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_15__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_5_15__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_16__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_16__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_17__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_17__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_18__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_18__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_19__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_19__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_20__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_20__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_21__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_21__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_22__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_22__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_23__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_5_23__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_24__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_24__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_25__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_25__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_26__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_26__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_27__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_27__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_28__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_28__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_29__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_29__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_30__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_30__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_5_31__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_5_31__leaf_clk));
 sky130_fd_sc_hd__inv_16 clkload0 (.A(clknet_5_0__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload1 (.A(clknet_5_1__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload2 (.A(clknet_5_2__leaf_clk));
 sky130_fd_sc_hd__inv_16 clkload3 (.A(clknet_5_3__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload4 (.A(clknet_5_4__leaf_clk));
 sky130_fd_sc_hd__inv_16 clkload5 (.A(clknet_5_6__leaf_clk));
 sky130_fd_sc_hd__inv_16 clkload6 (.A(clknet_5_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload7 (.A(clknet_5_10__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload8 (.A(clknet_5_11__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload9 (.A(clknet_5_13__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload10 (.A(clknet_5_14__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload11 (.A(clknet_5_15__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload12 (.A(clknet_5_17__leaf_clk));
 sky130_fd_sc_hd__clkinv_16 clkload13 (.A(clknet_5_18__leaf_clk));
 sky130_fd_sc_hd__inv_16 clkload14 (.A(clknet_5_19__leaf_clk));
 sky130_fd_sc_hd__inv_16 clkload15 (.A(clknet_5_20__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload16 (.A(clknet_5_21__leaf_clk));
 sky130_fd_sc_hd__clkinv_16 clkload17 (.A(clknet_5_22__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload18 (.A(clknet_5_23__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload19 (.A(clknet_5_24__leaf_clk));
 sky130_fd_sc_hd__clkinv_16 clkload20 (.A(clknet_5_25__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload21 (.A(clknet_5_27__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload22 (.A(clknet_5_28__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload23 (.A(clknet_5_29__leaf_clk));
 sky130_fd_sc_hd__clkinv_8 clkload24 (.A(clknet_5_30__leaf_clk));
 sky130_fd_sc_hd__clkinv_16 clkload25 (.A(clknet_5_31__leaf_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload26 (.A(clknet_leaf_273_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload27 (.A(clknet_leaf_274_clk));
 sky130_fd_sc_hd__clkinv_1 clkload28 (.A(clknet_leaf_283_clk));
 sky130_fd_sc_hd__bufinv_16 clkload29 (.A(clknet_leaf_284_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload30 (.A(clknet_leaf_285_clk));
 sky130_fd_sc_hd__clkinv_1 clkload31 (.A(clknet_leaf_286_clk));
 sky130_fd_sc_hd__clkinv_2 clkload32 (.A(clknet_leaf_288_clk));
 sky130_fd_sc_hd__inv_8 clkload33 (.A(clknet_leaf_289_clk));
 sky130_fd_sc_hd__bufinv_16 clkload34 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkinv_1 clkload35 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload36 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__bufinv_16 clkload37 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkinv_2 clkload38 (.A(clknet_leaf_278_clk));
 sky130_fd_sc_hd__inv_6 clkload39 (.A(clknet_leaf_279_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload40 (.A(clknet_leaf_281_clk));
 sky130_fd_sc_hd__bufinv_16 clkload41 (.A(clknet_leaf_282_clk));
 sky130_fd_sc_hd__bufinv_16 clkload42 (.A(clknet_leaf_287_clk));
 sky130_fd_sc_hd__inv_8 clkload43 (.A(clknet_leaf_290_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload44 (.A(clknet_leaf_263_clk));
 sky130_fd_sc_hd__clkinv_1 clkload45 (.A(clknet_leaf_264_clk));
 sky130_fd_sc_hd__clkinv_2 clkload46 (.A(clknet_leaf_265_clk));
 sky130_fd_sc_hd__clkinv_1 clkload47 (.A(clknet_leaf_266_clk));
 sky130_fd_sc_hd__clkinv_1 clkload48 (.A(clknet_leaf_267_clk));
 sky130_fd_sc_hd__bufinv_16 clkload49 (.A(clknet_leaf_268_clk));
 sky130_fd_sc_hd__clkinv_2 clkload50 (.A(clknet_leaf_269_clk));
 sky130_fd_sc_hd__clkinv_1 clkload51 (.A(clknet_leaf_270_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload52 (.A(clknet_leaf_275_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload53 (.A(clknet_leaf_256_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload54 (.A(clknet_leaf_257_clk));
 sky130_fd_sc_hd__clkinv_2 clkload55 (.A(clknet_leaf_259_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload56 (.A(clknet_leaf_260_clk));
 sky130_fd_sc_hd__clkinv_1 clkload57 (.A(clknet_leaf_261_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload58 (.A(clknet_leaf_276_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload59 (.A(clknet_leaf_277_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload60 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkinv_1 clkload61 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkinv_2 clkload62 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkinv_1 clkload63 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload64 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkinv_1 clkload65 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload66 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkinv_2 clkload67 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkinv_2 clkload68 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload69 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkinv_2 clkload70 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload71 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkinv_2 clkload72 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkinv_2 clkload73 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload74 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__bufinv_16 clkload75 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkinv_1 clkload76 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__bufinv_16 clkload77 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkinv_4 clkload78 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkinv_2 clkload79 (.A(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload80 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkinv_1 clkload81 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkinv_2 clkload82 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload83 (.A(clknet_leaf_248_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload84 (.A(clknet_leaf_251_clk));
 sky130_fd_sc_hd__clkinv_2 clkload85 (.A(clknet_leaf_252_clk));
 sky130_fd_sc_hd__clkinv_2 clkload86 (.A(clknet_leaf_253_clk));
 sky130_fd_sc_hd__bufinv_16 clkload87 (.A(clknet_leaf_254_clk));
 sky130_fd_sc_hd__clkinv_1 clkload88 (.A(clknet_leaf_255_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload89 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkinv_2 clkload90 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload91 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkinv_4 clkload92 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload93 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkinv_4 clkload94 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkinv_2 clkload95 (.A(clknet_leaf_38_clk));
 sky130_fd_sc_hd__inv_6 clkload96 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkinv_1 clkload97 (.A(clknet_leaf_218_clk));
 sky130_fd_sc_hd__bufinv_16 clkload98 (.A(clknet_leaf_219_clk));
 sky130_fd_sc_hd__clkinv_1 clkload99 (.A(clknet_leaf_220_clk));
 sky130_fd_sc_hd__clkinv_2 clkload100 (.A(clknet_leaf_221_clk));
 sky130_fd_sc_hd__bufinv_16 clkload101 (.A(clknet_leaf_222_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload102 (.A(clknet_leaf_223_clk));
 sky130_fd_sc_hd__clkinv_2 clkload103 (.A(clknet_leaf_224_clk));
 sky130_fd_sc_hd__bufinv_16 clkload104 (.A(clknet_leaf_225_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload105 (.A(clknet_leaf_226_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload106 (.A(clknet_leaf_228_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload107 (.A(clknet_leaf_229_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload108 (.A(clknet_leaf_230_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload109 (.A(clknet_leaf_231_clk));
 sky130_fd_sc_hd__clkinv_1 clkload110 (.A(clknet_leaf_234_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload111 (.A(clknet_leaf_235_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload112 (.A(clknet_leaf_238_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload113 (.A(clknet_leaf_239_clk));
 sky130_fd_sc_hd__clkinv_4 clkload114 (.A(clknet_leaf_209_clk));
 sky130_fd_sc_hd__clkinv_1 clkload115 (.A(clknet_leaf_210_clk));
 sky130_fd_sc_hd__inv_6 clkload116 (.A(clknet_leaf_211_clk));
 sky130_fd_sc_hd__clkinv_1 clkload117 (.A(clknet_leaf_212_clk));
 sky130_fd_sc_hd__bufinv_16 clkload118 (.A(clknet_leaf_213_clk));
 sky130_fd_sc_hd__clkinv_2 clkload119 (.A(clknet_leaf_214_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload120 (.A(clknet_leaf_215_clk));
 sky130_fd_sc_hd__bufinv_16 clkload121 (.A(clknet_leaf_216_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload122 (.A(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkinv_1 clkload123 (.A(clknet_leaf_202_clk));
 sky130_fd_sc_hd__clkinv_1 clkload124 (.A(clknet_leaf_203_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload125 (.A(clknet_leaf_205_clk));
 sky130_fd_sc_hd__clkinv_4 clkload126 (.A(clknet_leaf_206_clk));
 sky130_fd_sc_hd__bufinv_16 clkload127 (.A(clknet_leaf_207_clk));
 sky130_fd_sc_hd__bufinv_16 clkload128 (.A(clknet_leaf_217_clk));
 sky130_fd_sc_hd__bufinv_16 clkload129 (.A(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkinv_4 clkload130 (.A(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload131 (.A(clknet_leaf_237_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload132 (.A(clknet_leaf_240_clk));
 sky130_fd_sc_hd__clkbuf_16 clkload133 (.A(clknet_leaf_241_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload134 (.A(clknet_leaf_242_clk));
 sky130_fd_sc_hd__inv_4 clkload135 (.A(clknet_leaf_243_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload136 (.A(clknet_leaf_249_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload137 (.A(clknet_leaf_250_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload138 (.A(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload139 (.A(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload140 (.A(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkinv_1 clkload141 (.A(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload142 (.A(clknet_leaf_246_clk));
 sky130_fd_sc_hd__clkinv_2 clkload143 (.A(clknet_leaf_247_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload144 (.A(clknet_leaf_186_clk));
 sky130_fd_sc_hd__inv_6 clkload145 (.A(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload146 (.A(clknet_leaf_189_clk));
 sky130_fd_sc_hd__bufinv_16 clkload147 (.A(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload148 (.A(clknet_leaf_198_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload149 (.A(clknet_leaf_199_clk));
 sky130_fd_sc_hd__inv_6 clkload150 (.A(clknet_leaf_204_clk));
 sky130_fd_sc_hd__clkinv_1 clkload151 (.A(clknet_leaf_183_clk));
 sky130_fd_sc_hd__bufinv_16 clkload152 (.A(clknet_leaf_190_clk));
 sky130_fd_sc_hd__bufinv_16 clkload153 (.A(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload154 (.A(clknet_leaf_193_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload155 (.A(clknet_leaf_194_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload156 (.A(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload157 (.A(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkinv_2 clkload158 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload159 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__bufinv_16 clkload160 (.A(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload161 (.A(clknet_leaf_53_clk));
 sky130_fd_sc_hd__inv_6 clkload162 (.A(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkinv_1 clkload163 (.A(clknet_leaf_55_clk));
 sky130_fd_sc_hd__bufinv_16 clkload164 (.A(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload165 (.A(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkinv_4 clkload166 (.A(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkinv_2 clkload167 (.A(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkinv_2 clkload168 (.A(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload169 (.A(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload170 (.A(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkinv_1 clkload171 (.A(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload172 (.A(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload173 (.A(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkinv_1 clkload174 (.A(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload175 (.A(clknet_leaf_73_clk));
 sky130_fd_sc_hd__bufinv_16 clkload176 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload177 (.A(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload178 (.A(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkinv_2 clkload179 (.A(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload180 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload181 (.A(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload182 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkinv_1 clkload183 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkinv_1 clkload184 (.A(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkinv_2 clkload185 (.A(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkinv_1 clkload186 (.A(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkinv_2 clkload187 (.A(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkinv_1 clkload188 (.A(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkinv_2 clkload189 (.A(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkinv_1 clkload190 (.A(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload191 (.A(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkinv_2 clkload192 (.A(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkinv_1 clkload193 (.A(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkinv_4 clkload194 (.A(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload195 (.A(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkinv_2 clkload196 (.A(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload197 (.A(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkinv_1 clkload198 (.A(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkinv_1 clkload199 (.A(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkinv_1 clkload200 (.A(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkinv_1 clkload201 (.A(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload202 (.A(clknet_leaf_88_clk));
 sky130_fd_sc_hd__bufinv_16 clkload203 (.A(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkinv_2 clkload204 (.A(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload205 (.A(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload206 (.A(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload207 (.A(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkinv_1 clkload208 (.A(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkinv_2 clkload209 (.A(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkinv_1 clkload210 (.A(clknet_leaf_95_clk));
 sky130_fd_sc_hd__bufinv_16 clkload211 (.A(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkinv_1 clkload212 (.A(clknet_leaf_97_clk));
 sky130_fd_sc_hd__bufinv_16 clkload213 (.A(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkinv_1 clkload214 (.A(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkinv_1 clkload215 (.A(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkinv_2 clkload216 (.A(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkinv_2 clkload217 (.A(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkinv_1 clkload218 (.A(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload219 (.A(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload220 (.A(clknet_leaf_173_clk));
 sky130_fd_sc_hd__bufinv_16 clkload221 (.A(clknet_leaf_176_clk));
 sky130_fd_sc_hd__bufinv_16 clkload222 (.A(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkinv_2 clkload223 (.A(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkinv_2 clkload224 (.A(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload225 (.A(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkinv_1 clkload226 (.A(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload227 (.A(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkinv_1 clkload228 (.A(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkinv_2 clkload229 (.A(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload230 (.A(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkinv_1 clkload231 (.A(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkinv_1 clkload232 (.A(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload233 (.A(clknet_leaf_169_clk));
 sky130_fd_sc_hd__bufinv_16 clkload234 (.A(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkinv_4 clkload235 (.A(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload236 (.A(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkinv_4 clkload237 (.A(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkinv_2 clkload238 (.A(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkinv_4 clkload239 (.A(clknet_leaf_158_clk));
 sky130_fd_sc_hd__bufinv_16 clkload240 (.A(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload241 (.A(clknet_leaf_160_clk));
 sky130_fd_sc_hd__inv_6 clkload242 (.A(clknet_leaf_161_clk));
 sky130_fd_sc_hd__inv_6 clkload243 (.A(clknet_leaf_174_clk));
 sky130_fd_sc_hd__bufinv_16 clkload244 (.A(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkinv_2 clkload245 (.A(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkinv_2 clkload246 (.A(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload247 (.A(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkinv_2 clkload248 (.A(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload249 (.A(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload250 (.A(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload251 (.A(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload252 (.A(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload253 (.A(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkinv_1 clkload254 (.A(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload255 (.A(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload256 (.A(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkinv_1 clkload257 (.A(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkinv_2 clkload258 (.A(clknet_leaf_134_clk));
 sky130_fd_sc_hd__bufinv_16 clkload259 (.A(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload260 (.A(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_1 clkload261 (.A(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload262 (.A(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkinv_4 clkload263 (.A(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload264 (.A(clknet_leaf_153_clk));
 sky130_fd_sc_hd__buf_2 rebuffer1 (.A(\hash.CA1.S1.X[30] ),
    .X(net1040));
 sky130_fd_sc_hd__buf_2 rebuffer2 (.A(net1040),
    .X(net1041));
 sky130_fd_sc_hd__buf_2 rebuffer3 (.A(net1040),
    .X(net1042));
 sky130_fd_sc_hd__buf_2 rebuffer4 (.A(_06727_),
    .X(net1043));
 sky130_fd_sc_hd__buf_2 rebuffer5 (.A(_04475_),
    .X(net1044));
 sky130_fd_sc_hd__buf_2 rebuffer6 (.A(net1044),
    .X(net1045));
 sky130_fd_sc_hd__buf_2 rebuffer7 (.A(net1045),
    .X(net1046));
 sky130_fd_sc_hd__buf_2 rebuffer8 (.A(net1045),
    .X(net1047));
 sky130_fd_sc_hd__buf_2 rebuffer9 (.A(net1047),
    .X(net1048));
 sky130_fd_sc_hd__buf_6 rebuffer10 (.A(\hash.CA1.S0.X[25] ),
    .X(net1049));
 sky130_fd_sc_hd__buf_2 rebuffer11 (.A(_13330_),
    .X(net1050));
 sky130_fd_sc_hd__buf_6 rebuffer12 (.A(_04710_),
    .X(net1051));
 sky130_fd_sc_hd__buf_2 rebuffer13 (.A(_04509_),
    .X(net1052));
 sky130_fd_sc_hd__buf_6 rebuffer14 (.A(_04635_),
    .X(net1053));
 sky130_fd_sc_hd__nor2_2 clone15 (.A(net1055),
    .B(net344),
    .Y(net1054));
 sky130_fd_sc_hd__buf_2 rebuffer16 (.A(_06682_),
    .X(net1055));
 sky130_fd_sc_hd__buf_2 rebuffer17 (.A(_06689_),
    .X(net1056));
 sky130_fd_sc_hd__buf_2 rebuffer18 (.A(net1056),
    .X(net1057));
 sky130_fd_sc_hd__buf_2 rebuffer19 (.A(net1056),
    .X(net1058));
 sky130_fd_sc_hd__buf_2 rebuffer20 (.A(_13461_),
    .X(net1059));
 sky130_fd_sc_hd__buf_2 rebuffer21 (.A(\hash.CA2.S1.X[25] ),
    .X(net1060));
 sky130_fd_sc_hd__buf_2 rebuffer22 (.A(\hash.CA2.S1.X[25] ),
    .X(net1061));
 sky130_fd_sc_hd__buf_2 rebuffer23 (.A(\hash.CA2.S1.X[25] ),
    .X(net1062));
 sky130_fd_sc_hd__buf_2 rebuffer24 (.A(net1122),
    .X(net1063));
 sky130_fd_sc_hd__buf_2 rebuffer25 (.A(_13414_),
    .X(net1064));
 sky130_fd_sc_hd__buf_2 rebuffer26 (.A(_13351_),
    .X(net1065));
 sky130_fd_sc_hd__buf_6 rebuffer27 (.A(_13386_),
    .X(net1066));
 sky130_fd_sc_hd__buf_2 rebuffer28 (.A(net1066),
    .X(net1067));
 sky130_fd_sc_hd__buf_2 rebuffer29 (.A(_13379_),
    .X(net1068));
 sky130_fd_sc_hd__buf_2 rebuffer30 (.A(_04537_),
    .X(net1069));
 sky130_fd_sc_hd__buf_2 rebuffer31 (.A(net1069),
    .X(net1070));
 sky130_fd_sc_hd__buf_2 rebuffer32 (.A(net1069),
    .X(net1071));
 sky130_fd_sc_hd__buf_2 rebuffer33 (.A(_04537_),
    .X(net1072));
 sky130_fd_sc_hd__buf_2 rebuffer34 (.A(net1072),
    .X(net1073));
 sky130_fd_sc_hd__buf_2 rebuffer35 (.A(\hash.CA2.S1.X[6] ),
    .X(net1074));
 sky130_fd_sc_hd__buf_2 rebuffer36 (.A(\hash.CA2.S1.X[6] ),
    .X(net1075));
 sky130_fd_sc_hd__buf_2 rebuffer37 (.A(net1075),
    .X(net1076));
 sky130_fd_sc_hd__buf_2 rebuffer38 (.A(net1076),
    .X(net1077));
 sky130_fd_sc_hd__buf_2 rebuffer39 (.A(_04612_),
    .X(net1078));
 sky130_fd_sc_hd__buf_2 rebuffer40 (.A(net1078),
    .X(net1079));
 sky130_fd_sc_hd__buf_2 rebuffer41 (.A(\hash.CA2.S1.X[7] ),
    .X(net1080));
 sky130_fd_sc_hd__buf_2 rebuffer42 (.A(\hash.CA2.S1.X[7] ),
    .X(net1081));
 sky130_fd_sc_hd__buf_2 rebuffer43 (.A(net1081),
    .X(net1082));
 sky130_fd_sc_hd__buf_2 rebuffer44 (.A(net1081),
    .X(net1083));
 sky130_fd_sc_hd__buf_2 rebuffer45 (.A(net1081),
    .X(net1084));
 sky130_fd_sc_hd__buf_2 rebuffer46 (.A(_04402_),
    .X(net1085));
 sky130_fd_sc_hd__buf_2 rebuffer47 (.A(\hash.CA2.S1.X[26] ),
    .X(net1086));
 sky130_fd_sc_hd__buf_2 rebuffer48 (.A(\hash.CA2.S1.X[26] ),
    .X(net1087));
 sky130_fd_sc_hd__buf_2 rebuffer49 (.A(_12086_),
    .X(net1088));
 sky130_fd_sc_hd__buf_2 rebuffer50 (.A(_13237_),
    .X(net1089));
 sky130_fd_sc_hd__buf_2 rebuffer51 (.A(_04688_),
    .X(net1090));
 sky130_fd_sc_hd__buf_2 rebuffer52 (.A(_06151_),
    .X(net1091));
 sky130_fd_sc_hd__buf_2 rebuffer53 (.A(\hash.CA2.S1.X[25] ),
    .X(net1092));
 sky130_fd_sc_hd__buf_2 rebuffer60 (.A(_13344_),
    .X(net1099));
 sky130_fd_sc_hd__buf_2 rebuffer61 (.A(\hash.CA2.S1.X[26] ),
    .X(net1100));
 sky130_fd_sc_hd__buf_2 rebuffer68 (.A(_04481_),
    .X(net1107));
 sky130_fd_sc_hd__buf_2 rebuffer69 (.A(_06045_),
    .X(net1108));
 sky130_fd_sc_hd__buf_2 rebuffer72 (.A(_09231_),
    .X(net1111));
 sky130_fd_sc_hd__mux2i_4 clone73 (.A0(\w[63][24] ),
    .A1(_05325_),
    .S(net339),
    .Y(net1112));
 sky130_fd_sc_hd__a21oi_4 clone74 (.A1(\w[63][28] ),
    .A2(done),
    .B1(_05371_),
    .Y(net1113));
 sky130_fd_sc_hd__a21oi_4 clone75 (.A1(\w[63][30] ),
    .A2(net355),
    .B1(_05388_),
    .Y(net1114));
 sky130_fd_sc_hd__buf_8 load_slew1 (.A(\count2_1[1] ),
    .X(net1093));
 sky130_fd_sc_hd__buf_2 rebuffer15 (.A(_06952_),
    .X(net1094));
 sky130_fd_sc_hd__buf_12 rebuffer54 (.A(_04588_),
    .X(net1095));
 sky130_fd_sc_hd__buf_2 rebuffer55 (.A(_04472_),
    .X(net1096));
 sky130_fd_sc_hd__o22a_2 clone56 (.A1(net345),
    .A2(_06705_),
    .B1(_06706_),
    .B2(_06704_),
    .X(net1097));
 sky130_fd_sc_hd__buf_2 rebuffer57 (.A(_12728_),
    .X(net1098));
 sky130_fd_sc_hd__buf_2 rebuffer58 (.A(_04517_),
    .X(net1101));
 sky130_fd_sc_hd__buf_2 rebuffer59 (.A(net1101),
    .X(net1102));
 sky130_fd_sc_hd__buf_2 rebuffer62 (.A(net1101),
    .X(net1103));
 sky130_fd_sc_hd__buf_2 rebuffer63 (.A(\hash.CA2.S1.X[1] ),
    .X(net1104));
 sky130_fd_sc_hd__buf_2 rebuffer64 (.A(\hash.CA2.S1.X[1] ),
    .X(net1105));
 sky130_fd_sc_hd__buf_4 rebuffer67 (.A(\hash.CA2.S1.X[8] ),
    .X(net1110));
 sky130_fd_sc_hd__buf_2 rebuffer70 (.A(\hash.CA2.S1.X[8] ),
    .X(net1115));
 sky130_fd_sc_hd__buf_2 rebuffer71 (.A(net1115),
    .X(net1116));
 sky130_fd_sc_hd__buf_2 rebuffer73 (.A(net1116),
    .X(net1117));
 sky130_fd_sc_hd__buf_2 rebuffer74 (.A(\hash.CA2.S1.X[27] ),
    .X(net1118));
 sky130_fd_sc_hd__buf_2 rebuffer75 (.A(\hash.CA2.S1.X[2] ),
    .X(net1119));
 sky130_fd_sc_hd__buf_2 rebuffer76 (.A(net1119),
    .X(net1120));
 sky130_fd_sc_hd__buf_2 rebuffer77 (.A(\hash.CA2.S1.X[2] ),
    .X(net1121));
 sky130_fd_sc_hd__buf_2 rebuffer78 (.A(\hash.CA2.S1.X[25] ),
    .X(net1122));
 sky130_fd_sc_hd__buf_6 rebuffer79 (.A(_06710_),
    .X(net1123));
 sky130_fd_sc_hd__buf_2 rebuffer80 (.A(_06699_),
    .X(net1124));
 sky130_fd_sc_hd__buf_2 rebuffer81 (.A(_13245_),
    .X(net1125));
 sky130_fd_sc_hd__buf_12 rebuffer83 (.A(_06164_),
    .X(net1127));
 sky130_fd_sc_hd__a21oi_4 clone84 (.A1(\w[62][24] ),
    .A2(net353),
    .B1(_04999_),
    .Y(net1128));
 sky130_fd_sc_hd__buf_12 rebuffer85 (.A(_05000_),
    .X(net1129));
 sky130_fd_sc_hd__clkbuf_4 split89 (.A(\count15_2[2] ),
    .X(net1133));
 sky130_fd_sc_hd__a21oi_2 clone90 (.A1(\w[63][28] ),
    .A2(done),
    .B1(_05371_),
    .Y(net1134));
 sky130_fd_sc_hd__mux2i_4 clone91 (.A0(\w[62][28] ),
    .A1(_05034_),
    .S(_04797_),
    .Y(net1135));
 sky130_fd_sc_hd__a21oi_4 clone92 (.A1(\w[63][18] ),
    .A2(net350),
    .B1(_05266_),
    .Y(net1136));
 sky130_fd_sc_hd__a21oi_2 clone93 (.A1(\w[62][22] ),
    .A2(net353),
    .B1(_04983_),
    .Y(net1137));
 sky130_fd_sc_hd__a21oi_4 clone94 (.A1(\w[63][14] ),
    .A2(net350),
    .B1(_05227_),
    .Y(net1138));
 sky130_fd_sc_hd__a21oi_4 clone95 (.A1(\w[62][26] ),
    .A2(net353),
    .B1(_05019_),
    .Y(net1139));
 sky130_fd_sc_hd__a21oi_4 clone96 (.A1(\w[63][16] ),
    .A2(net351),
    .B1(_05246_),
    .Y(net1140));
 sky130_fd_sc_hd__a21oi_2 clone97 (.A1(\w[63][28] ),
    .A2(done),
    .B1(_05371_),
    .Y(net1141));
 sky130_fd_sc_hd__a21oi_2 clone98 (.A1(\w[62][18] ),
    .A2(net352),
    .B1(_04938_),
    .Y(net1142));
 sky130_fd_sc_hd__buf_12 rebuffer99 (.A(_05389_),
    .X(net1143));
 sky130_fd_sc_hd__o21ai_2 clone100 (.A1(\w[63][26] ),
    .A2(net339),
    .B1(_05346_),
    .Y(net1144));
 sky130_fd_sc_hd__buf_12 rebuffer101 (.A(_05326_),
    .X(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_00006_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_00008_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_00017_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_00017_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_00017_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(_00024_));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(_00024_));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(_00024_));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(_00024_));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(_00024_));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(_00024_));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(_00025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(_00026_));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(_00029_));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(_00052_));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(_00055_));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(_00058_));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(_00061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(_00061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(_00061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(_00061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(_00061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(_00061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(_00061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(_00061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(_00061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(_00061_));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(_00063_));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(_00063_));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(_00063_));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(_00063_));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(_00063_));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(_00063_));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(_00063_));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(_00092_));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(_09009_));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(_09130_));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(_11620_));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(_11748_));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(_11756_));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(_11979_));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(_12019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(\hash.CA1.p3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(\hash.CA1.p3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(\hash.CA1.p3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(\hash.CA1.p3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(\hash.CA1.p3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(\hash.CA1.p3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(\hash.CA1.p3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(\hash.CA1.p3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(\hash.CA1.p3[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(\hash.CA1.p3[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(\hash.CA1.p3[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(\hash.CA1.p3[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(\hash.CA1.p3[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(_00028_));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(_00050_));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(_00021_));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(_00023_));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(_00020_));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(_00002_));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(_00019_));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(_00039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(_00040_));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(_00043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(_00043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(_00043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(_00043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(_00043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(_00047_));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(_00047_));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(_00047_));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(_00047_));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(_00047_));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(_00051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(_00126_));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(_06747_));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(_08960_));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(_09150_));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(_11586_));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(_12368_));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(\hash.CA1.S1.X[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(\hash.CA1.S1.X[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(\hash.CA1.p2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(net854));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(_00007_));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(_00047_));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(_00047_));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(_00051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(_00051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(_00051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(\hash.CA1.p2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(_00051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(_00051_));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(\hash.CA1.p2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(\hash.CA1.p2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(\hash.CA1.p2[0] ));
 sky130_fd_sc_hd__fill_8 FILLER_0_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_374 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_536 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_680 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_788 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_817 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1427 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1457 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_0_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_0_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_558 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_574 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_754 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_908 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_983 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_990 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_998 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_1_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_1_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_952 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_2_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_2_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_636 ();
 sky130_fd_sc_hd__fill_4 FILLER_3_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_3_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_830 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_4_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_4_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_400 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_696 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_5_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_826 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_5_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_393 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_6_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_6_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_267 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_450 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_855 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_7_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_7_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_845 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_8_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_8_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_493 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_9_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_9_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_657 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_744 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_10_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_10_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_321 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_11_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_876 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_11_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_315 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_12_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_12_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_284 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_844 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_13_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_13_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_14_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_14_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_512 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_15_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_15_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_422 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_16_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_16_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_520 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_17_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_870 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_17_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_704 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_934 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_950 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_966 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_18_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_18_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_270 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_813 ();
 sky130_fd_sc_hd__fill_4 FILLER_19_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_19_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_771 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_20_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_20_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_552 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_604 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_21_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1353 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_21_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_177 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_297 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_484 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_960 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1286 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_22_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_22_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_201 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_406 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_604 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_692 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_913 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_938 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1235 ();
 sky130_fd_sc_hd__fill_4 FILLER_23_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1267 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1280 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_23_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_537 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1205 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1226 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1262 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1270 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1325 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1355 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_24_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_24_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1236 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1287 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1312 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1365 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1427 ();
 sky130_fd_sc_hd__fill_4 FILLER_25_1435 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_25_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_480 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_768 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_829 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1300 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1326 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1382 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1390 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1398 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_1406 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1435 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1445 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_26_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_26_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1188 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1209 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1223 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1325 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_27_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1404 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_27_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_713 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1294 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1302 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1310 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1314 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1338 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1342 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1359 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_28_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_28_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_930 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1040 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1206 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1214 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1258 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1316 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1366 ();
 sky130_fd_sc_hd__fill_4 FILLER_29_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_29_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_773 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_835 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1273 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1295 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1301 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1419 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1427 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1450 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1458 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1466 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_30_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_30_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_501 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_927 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1172 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1233 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1272 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1281 ();
 sky130_fd_sc_hd__fill_4 FILLER_31_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1312 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1354 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1439 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1466 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1474 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1482 ();
 sky130_fd_sc_hd__fill_8 FILLER_31_1490 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_374 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_660 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_720 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1082 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1178 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1200 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1303 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1376 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1384 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1392 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1400 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1408 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1452 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1460 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1468 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_32_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_32_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_210 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_276 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_606 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_863 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_873 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_934 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1103 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1232 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1285 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1304 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1347 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1370 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1376 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1430 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1438 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1468 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1476 ();
 sky130_fd_sc_hd__fill_8 FILLER_33_1484 ();
 sky130_fd_sc_hd__fill_4 FILLER_33_1492 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1496 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_368 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_534 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_829 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1099 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1320 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1359 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1403 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1409 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1434 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1438 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1464 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1468 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_34_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_34_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_512 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_550 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_608 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_612 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_987 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1123 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1256 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1303 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1316 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1340 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1346 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1350 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1360 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1398 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1403 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1407 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1424 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1432 ();
 sky130_fd_sc_hd__fill_4 FILLER_35_1436 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1448 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1456 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1464 ();
 sky130_fd_sc_hd__fill_8 FILLER_35_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_773 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1099 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1159 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1233 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1309 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1318 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1320 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1358 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1375 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1409 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1434 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1453 ();
 sky130_fd_sc_hd__fill_8 FILLER_36_1461 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1469 ();
 sky130_fd_sc_hd__fill_4 FILLER_36_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_831 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_892 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_984 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_992 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1000 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1103 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1170 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1223 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1265 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1308 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1316 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1335 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1347 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1363 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1390 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1392 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1400 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1425 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1438 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_37_1486 ();
 sky130_fd_sc_hd__fill_4 FILLER_37_1494 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_182 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1015 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1207 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1226 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1357 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1377 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1423 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1452 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1460 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1468 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1477 ();
 sky130_fd_sc_hd__fill_8 FILLER_38_1485 ();
 sky130_fd_sc_hd__fill_4 FILLER_38_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_913 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1083 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1369 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1388 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1396 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1404 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1412 ();
 sky130_fd_sc_hd__fill_4 FILLER_39_1436 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_39_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_463 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_502 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_522 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_782 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_897 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1077 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1257 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1267 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1361 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1375 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1431 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1474 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1478 ();
 sky130_fd_sc_hd__fill_8 FILLER_40_1486 ();
 sky130_fd_sc_hd__fill_4 FILLER_40_1494 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_200 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_452 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_990 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_998 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1224 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1242 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_41_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_41_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1494 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_550 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_953 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1238 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1249 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1270 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1298 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1306 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1314 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_42_1377 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1409 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1425 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1427 ();
 sky130_fd_sc_hd__fill_4 FILLER_42_1445 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_184 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_332 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1105 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1136 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1183 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1216 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1333 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1366 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1371 ();
 sky130_fd_sc_hd__fill_4 FILLER_43_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1406 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1414 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1422 ();
 sky130_fd_sc_hd__fill_8 FILLER_43_1430 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1438 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1472 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_420 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_837 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1014 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1022 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1077 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1114 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1304 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1327 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1338 ();
 sky130_fd_sc_hd__fill_4 FILLER_44_1346 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1372 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1393 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_44_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1459 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1461 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1161 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1220 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1271 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1281 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1292 ();
 sky130_fd_sc_hd__fill_8 FILLER_45_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1355 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1376 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1404 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1408 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1433 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1439 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1473 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1490 ();
 sky130_fd_sc_hd__fill_4 FILLER_45_1494 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_351 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_594 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_852 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1015 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1058 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1070 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1088 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1135 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1160 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1270 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1364 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1372 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1376 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1378 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1386 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1400 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1408 ();
 sky130_fd_sc_hd__fill_8 FILLER_46_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1446 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1464 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1468 ();
 sky130_fd_sc_hd__fill_4 FILLER_46_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1087 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1095 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1110 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1122 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1213 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1287 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1327 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1388 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1400 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1408 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1412 ();
 sky130_fd_sc_hd__fill_4 FILLER_47_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_47_1464 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1472 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1474 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_300 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_590 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_606 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_620 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1014 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1022 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1030 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1044 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1094 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1134 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1288 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1305 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1313 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1364 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1372 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1380 ();
 sky130_fd_sc_hd__fill_8 FILLER_48_1400 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1408 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1438 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1440 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1454 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1458 ();
 sky130_fd_sc_hd__fill_4 FILLER_48_1466 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1471 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_522 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_618 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_801 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_970 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_978 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1054 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1095 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1177 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1240 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1286 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1298 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1313 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1325 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1338 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1342 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1357 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1365 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1369 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1441 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1449 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1453 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1455 ();
 sky130_fd_sc_hd__fill_8 FILLER_49_1464 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1472 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1476 ();
 sky130_fd_sc_hd__fill_4 FILLER_49_1483 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1487 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1494 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_364 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_758 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_970 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1023 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1100 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1288 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1323 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1362 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1370 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1396 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1398 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1406 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1417 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1434 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1442 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1446 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1463 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_50_1477 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_50_1491 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_516 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_670 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1116 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1167 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1175 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1227 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1302 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1335 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1365 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1395 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1403 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1407 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1421 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1433 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1439 ();
 sky130_fd_sc_hd__fill_4 FILLER_51_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_51_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_600 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_717 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_910 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_978 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1086 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1152 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1205 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1315 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1325 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1375 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1408 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1433 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_52_1474 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1482 ();
 sky130_fd_sc_hd__fill_4 FILLER_52_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1496 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_730 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_919 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_994 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1120 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1163 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1176 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1308 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1334 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1342 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1350 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1354 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1366 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1392 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1394 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1435 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1439 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_53_1481 ();
 sky130_fd_sc_hd__fill_4 FILLER_53_1492 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_662 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_938 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1118 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1313 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1318 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1330 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1336 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1368 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1384 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1386 ();
 sky130_fd_sc_hd__fill_8 FILLER_54_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1425 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1427 ();
 sky130_fd_sc_hd__fill_4 FILLER_54_1432 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1436 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1438 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_576 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_770 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_880 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1045 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1107 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1227 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1275 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1283 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1306 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1318 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1332 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1340 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1346 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1354 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1358 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1412 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1420 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1428 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1436 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1445 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1453 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1464 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1466 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1470 ();
 sky130_fd_sc_hd__fill_8 FILLER_55_1478 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1486 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1490 ();
 sky130_fd_sc_hd__fill_4 FILLER_55_1494 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_250 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_717 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_893 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_966 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_982 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1152 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1213 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1262 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1270 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1278 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1286 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1403 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1409 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1440 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1448 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_56_1479 ();
 sky130_fd_sc_hd__fill_4 FILLER_56_1487 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1491 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_252 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_452 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_507 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_570 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_903 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1120 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1128 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1136 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1161 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1304 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1312 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1329 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1410 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1412 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1432 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1434 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1438 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1441 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1449 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1459 ();
 sky130_fd_sc_hd__fill_8 FILLER_57_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1479 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1487 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1489 ();
 sky130_fd_sc_hd__fill_4 FILLER_57_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_971 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1210 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1235 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1308 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1324 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1332 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1402 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1420 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1428 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1432 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1450 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1452 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1460 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1462 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1468 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1474 ();
 sky130_fd_sc_hd__fill_4 FILLER_58_1482 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1486 ();
 sky130_fd_sc_hd__fill_8 FILLER_58_1490 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_138 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_270 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_828 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_907 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_971 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_990 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1223 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1244 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1253 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1329 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1388 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1417 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1425 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1433 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1439 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1445 ();
 sky130_fd_sc_hd__fill_4 FILLER_59_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1455 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1475 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1483 ();
 sky130_fd_sc_hd__fill_8 FILLER_59_1491 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_604 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1128 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1189 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1260 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1264 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1279 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1320 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1400 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1435 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1445 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_60_1479 ();
 sky130_fd_sc_hd__fill_4 FILLER_60_1487 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1491 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_804 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1052 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1107 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1176 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1222 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1283 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1287 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1387 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1395 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1403 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_61_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1445 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1455 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_61_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_111 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_187 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_775 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1073 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1080 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1116 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1148 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1193 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1331 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1339 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1357 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1384 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1392 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1400 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1408 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1447 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1453 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1468 ();
 sky130_fd_sc_hd__fill_8 FILLER_62_1484 ();
 sky130_fd_sc_hd__fill_4 FILLER_62_1492 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1496 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_204 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_512 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_700 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1056 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1123 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1174 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1304 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1312 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1348 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1356 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1358 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1366 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1401 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1409 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1417 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1459 ();
 sky130_fd_sc_hd__fill_8 FILLER_63_1467 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1475 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1482 ();
 sky130_fd_sc_hd__fill_4 FILLER_63_1491 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_288 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_378 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_540 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_724 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_815 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1057 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1069 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1205 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1257 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1272 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1288 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1314 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1326 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1334 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1346 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1376 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1423 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1444 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1446 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1453 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1464 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1468 ();
 sky130_fd_sc_hd__fill_8 FILLER_64_1471 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1479 ();
 sky130_fd_sc_hd__fill_4 FILLER_64_1486 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1490 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1492 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_469 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_555 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1054 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1087 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1101 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1223 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1312 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_65_1353 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1365 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1402 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1413 ();
 sky130_fd_sc_hd__fill_4 FILLER_65_1427 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_717 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_782 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_834 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1023 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1125 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1133 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1173 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1308 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1324 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1332 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1334 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1346 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1395 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1406 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1435 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1445 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1449 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1453 ();
 sky130_fd_sc_hd__fill_8 FILLER_66_1458 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1466 ();
 sky130_fd_sc_hd__fill_4 FILLER_66_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_383 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_966 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1091 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1122 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1281 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1305 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1327 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1338 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1346 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1350 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1362 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1423 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1441 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1449 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1453 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1455 ();
 sky130_fd_sc_hd__fill_8 FILLER_67_1472 ();
 sky130_fd_sc_hd__fill_4 FILLER_67_1480 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1484 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1486 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_132 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_220 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_386 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_474 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_482 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1020 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1104 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1114 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1286 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1362 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1374 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1395 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1420 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1422 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1426 ();
 sky130_fd_sc_hd__fill_8 FILLER_68_1434 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1453 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1474 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1476 ();
 sky130_fd_sc_hd__fill_4 FILLER_68_1480 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1484 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1491 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_127 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1091 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1150 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1279 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1287 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1302 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1372 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1412 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1428 ();
 sky130_fd_sc_hd__fill_4 FILLER_69_1436 ();
 sky130_fd_sc_hd__fill_8 FILLER_69_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_668 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_726 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_771 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1093 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1101 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1210 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1226 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1235 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1306 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1338 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1340 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1408 ();
 sky130_fd_sc_hd__fill_8 FILLER_70_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_70_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1445 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1473 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_95 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_200 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_593 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_607 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_817 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_893 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1101 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1151 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1203 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1239 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1273 ();
 sky130_fd_sc_hd__fill_4 FILLER_71_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1338 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1346 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1364 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1372 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_71_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1465 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_89 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_97 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_406 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_434 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_766 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1070 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1080 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1131 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1257 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1270 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1278 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1286 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1298 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1306 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1317 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1414 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1416 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1426 ();
 sky130_fd_sc_hd__fill_8 FILLER_72_1434 ();
 sky130_fd_sc_hd__fill_4 FILLER_72_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1497 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_133 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_564 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_604 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_678 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_998 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1100 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1215 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1225 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1240 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1303 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1311 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1376 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_73_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1449 ();
 sky130_fd_sc_hd__fill_4 FILLER_73_1458 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1462 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1464 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1497 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_18 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_533 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_790 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1032 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1077 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1190 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1202 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1233 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1253 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1310 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1324 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1333 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1369 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1394 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1402 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1406 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1419 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1425 ();
 sky130_fd_sc_hd__fill_4 FILLER_74_1433 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1444 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1452 ();
 sky130_fd_sc_hd__fill_8 FILLER_74_1460 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1468 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1471 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1497 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_118 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_135 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_995 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1023 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1033 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1101 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1120 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1339 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1343 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1360 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1393 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1409 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1413 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1430 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1434 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_75_1457 ();
 sky130_fd_sc_hd__fill_4 FILLER_75_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_63 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_950 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1028 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1082 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1129 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1182 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1209 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1251 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1266 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1296 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1323 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1325 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1338 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1346 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1361 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1375 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1436 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1445 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_76_1476 ();
 sky130_fd_sc_hd__fill_4 FILLER_76_1484 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1488 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_90 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_98 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_198 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_263 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_418 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_576 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1304 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1312 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1342 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1372 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1398 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1400 ();
 sky130_fd_sc_hd__fill_4 FILLER_77_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1430 ();
 sky130_fd_sc_hd__fill_8 FILLER_77_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_117 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_218 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_604 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_782 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1134 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1215 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1254 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1262 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1271 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_78_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1431 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_78_1487 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1495 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_305 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_847 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_878 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1061 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1086 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1104 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1240 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1298 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1368 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1376 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1398 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1406 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1410 ();
 sky130_fd_sc_hd__fill_8 FILLER_79_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1424 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1445 ();
 sky130_fd_sc_hd__fill_4 FILLER_79_1462 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1466 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1468 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1496 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_910 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_952 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1125 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1173 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1204 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1258 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1267 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1273 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1333 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1359 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1372 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1387 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1396 ();
 sky130_fd_sc_hd__fill_4 FILLER_80_1404 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1408 ();
 sky130_fd_sc_hd__fill_8 FILLER_80_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1471 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1497 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_375 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_484 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_520 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_680 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_694 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_740 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_934 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1177 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1220 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1234 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1242 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1378 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1436 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1452 ();
 sky130_fd_sc_hd__fill_8 FILLER_81_1480 ();
 sky130_fd_sc_hd__fill_4 FILLER_81_1491 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_82 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_808 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_846 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_862 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_904 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1098 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1102 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1135 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1298 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1306 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1314 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1322 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1330 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1338 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1346 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1364 ();
 sky130_fd_sc_hd__fill_8 FILLER_82_1388 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1396 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1409 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1447 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1453 ();
 sky130_fd_sc_hd__fill_4 FILLER_82_1471 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_21 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_37 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_45 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_452 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_904 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1115 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1198 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1258 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1281 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1332 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1344 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1350 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1354 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1384 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1392 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1405 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_83_1432 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1462 ();
 sky130_fd_sc_hd__fill_4 FILLER_83_1488 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1492 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1496 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_88 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_105 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_130 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_936 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1190 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1260 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1332 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1372 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1374 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1457 ();
 sky130_fd_sc_hd__fill_4 FILLER_84_1465 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_84_1487 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1495 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_5 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_87 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_452 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_528 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_596 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_867 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_978 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1039 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1060 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1110 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1122 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1225 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1272 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1284 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1325 ();
 sky130_fd_sc_hd__fill_4 FILLER_85_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1401 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1432 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1452 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1458 ();
 sky130_fd_sc_hd__fill_8 FILLER_85_1463 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1473 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_426 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_724 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1015 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1140 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1161 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1222 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1240 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1248 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1256 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1264 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1326 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1334 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1342 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1393 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_86_1456 ();
 sky130_fd_sc_hd__fill_4 FILLER_86_1464 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1468 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1498 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_81 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_807 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1039 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1227 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1279 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1346 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1354 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1360 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1438 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1445 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1453 ();
 sky130_fd_sc_hd__fill_8 FILLER_87_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1465 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1467 ();
 sky130_fd_sc_hd__fill_4 FILLER_87_1492 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1496 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_302 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_420 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_723 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_784 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_822 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_880 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1189 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1251 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1369 ();
 sky130_fd_sc_hd__fill_8 FILLER_88_1384 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1426 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1428 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1445 ();
 sky130_fd_sc_hd__fill_4 FILLER_88_1463 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_366 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_580 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_732 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1050 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1061 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1102 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1156 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1164 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1172 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1225 ();
 sky130_fd_sc_hd__fill_4 FILLER_89_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1280 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1288 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1296 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1365 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1386 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1434 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1459 ();
 sky130_fd_sc_hd__fill_8 FILLER_89_1488 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_96 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_104 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_471 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_600 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_882 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1062 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1118 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1146 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1203 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1250 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1266 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1336 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1348 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1390 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1398 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1406 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1437 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1445 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1447 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_90_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1469 ();
 sky130_fd_sc_hd__fill_4 FILLER_90_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_94 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_102 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_156 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_203 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_327 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_402 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_874 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1162 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1170 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1280 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1288 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1296 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1327 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1343 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1347 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1396 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1404 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1418 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1433 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1439 ();
 sky130_fd_sc_hd__fill_4 FILLER_91_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_91_1461 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1469 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1473 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_357 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_405 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_645 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_964 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1262 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1270 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_92_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1323 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1335 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1418 ();
 sky130_fd_sc_hd__fill_4 FILLER_92_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1453 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1474 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_499 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_624 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1040 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1093 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1258 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1286 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1344 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1346 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1357 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1403 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1420 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1424 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1434 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1438 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1441 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1452 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1456 ();
 sky130_fd_sc_hd__fill_4 FILLER_93_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_93_1488 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_256 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_278 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_348 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_368 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_660 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_674 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1026 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1150 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1188 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1249 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1276 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1314 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1322 ();
 sky130_fd_sc_hd__fill_4 FILLER_94_1346 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1424 ();
 sky130_fd_sc_hd__fill_8 FILLER_94_1432 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1440 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1465 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_8 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_95 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_284 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_330 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1000 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1054 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1062 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1116 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1136 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1156 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1164 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1265 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1344 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1352 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1434 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1441 ();
 sky130_fd_sc_hd__fill_4 FILLER_95_1449 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1453 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_95_1487 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_542 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_714 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_806 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1034 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1061 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1245 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1253 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1313 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1391 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1403 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1409 ();
 sky130_fd_sc_hd__fill_4 FILLER_96_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1417 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1437 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1445 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1453 ();
 sky130_fd_sc_hd__fill_8 FILLER_96_1461 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_100 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_683 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_994 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1040 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1052 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1072 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1114 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1183 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1332 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1340 ();
 sky130_fd_sc_hd__fill_8 FILLER_97_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_97_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1398 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1445 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1450 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1458 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1487 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1493 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_900 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_995 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1077 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1142 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1152 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1214 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1251 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1268 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1364 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_98_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1469 ();
 sky130_fd_sc_hd__fill_4 FILLER_98_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_443 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_640 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_923 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_951 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_987 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1076 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1101 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1132 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1152 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1167 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1198 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1305 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1353 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1368 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1376 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1387 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1395 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1399 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1439 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1445 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1473 ();
 sky130_fd_sc_hd__fill_4 FILLER_99_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1485 ();
 sky130_fd_sc_hd__fill_8 FILLER_99_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_103 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_542 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_591 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_724 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_856 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_949 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_957 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1070 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1251 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1369 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1386 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1398 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1400 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1404 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1424 ();
 sky130_fd_sc_hd__fill_8 FILLER_100_1432 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1440 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1469 ();
 sky130_fd_sc_hd__fill_4 FILLER_100_1471 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_133 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_461 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_504 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_536 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_864 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1000 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1047 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1069 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1183 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1387 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1427 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1435 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1439 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_101_1472 ();
 sky130_fd_sc_hd__fill_4 FILLER_101_1480 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1487 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1493 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_354 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_577 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_606 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_666 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_980 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1022 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1077 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1123 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1142 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1197 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1267 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1275 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1375 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1425 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1433 ();
 sky130_fd_sc_hd__fill_4 FILLER_102_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1445 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1476 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1484 ();
 sky130_fd_sc_hd__fill_8 FILLER_102_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_85 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_192 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_218 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_443 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_506 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_564 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_765 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_952 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1100 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1131 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1136 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1159 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1167 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1175 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1339 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_103_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1441 ();
 sky130_fd_sc_hd__fill_4 FILLER_103_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1493 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1495 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_224 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_717 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1000 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1137 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1188 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1196 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1363 ();
 sky130_fd_sc_hd__fill_8 FILLER_104_1371 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1385 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1415 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1440 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1444 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1471 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1475 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1481 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1489 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1491 ();
 sky130_fd_sc_hd__fill_4 FILLER_104_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_69 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_92 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_143 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_821 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_963 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_992 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1086 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1120 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1189 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1219 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1282 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1290 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1292 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1338 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1358 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1366 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1378 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1423 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1427 ();
 sky130_fd_sc_hd__fill_4 FILLER_105_1435 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1439 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_105_1477 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1490 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1492 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_79 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_371 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_535 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_602 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_618 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_709 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_736 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_913 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1004 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1066 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1086 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1129 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1137 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1214 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1246 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1318 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1388 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1396 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1398 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1406 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_106_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_106_1495 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_10 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_694 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_741 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1002 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1014 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1240 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1310 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1312 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1342 ();
 sky130_fd_sc_hd__fill_4 FILLER_107_1350 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1354 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1379 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1422 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1480 ();
 sky130_fd_sc_hd__fill_8 FILLER_107_1488 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_474 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_518 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_722 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_954 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_981 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1073 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1197 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1205 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1238 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1302 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_108_1369 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1377 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1420 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1422 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1435 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1468 ();
 sky130_fd_sc_hd__fill_4 FILLER_108_1487 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1491 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_12 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_476 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_495 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_713 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_760 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_787 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_936 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_944 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_987 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1011 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1107 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1190 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1212 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1240 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1298 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1302 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1313 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_109_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1406 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1438 ();
 sky130_fd_sc_hd__fill_4 FILLER_109_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_83 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_97 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_537 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_840 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_893 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_968 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_985 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1011 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1016 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1020 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1083 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1101 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1237 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1376 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1378 ();
 sky130_fd_sc_hd__fill_4 FILLER_110_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1417 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1428 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_110_1479 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1487 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1489 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_118 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_160 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_484 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_501 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_553 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_709 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_945 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_976 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_996 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1015 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1062 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1107 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1232 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1250 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1278 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1288 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1390 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1398 ();
 sky130_fd_sc_hd__fill_4 FILLER_111_1406 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1410 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1412 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1465 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1476 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1478 ();
 sky130_fd_sc_hd__fill_8 FILLER_111_1482 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_148 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_177 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_240 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_277 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_372 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_443 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_470 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_540 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_738 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_874 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_912 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1010 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1263 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1275 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1315 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_112_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1427 ();
 sky130_fd_sc_hd__fill_4 FILLER_112_1466 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1495 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_674 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_728 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_892 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_972 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_980 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1046 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1226 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1295 ();
 sky130_fd_sc_hd__fill_4 FILLER_113_1316 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1366 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1439 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1448 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1450 ();
 sky130_fd_sc_hd__fill_8 FILLER_113_1454 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1462 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_71 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_650 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_787 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_900 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_908 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1023 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1040 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1069 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1077 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1393 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_114_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1419 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1423 ();
 sky130_fd_sc_hd__fill_4 FILLER_114_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1445 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_79 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_580 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_810 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_895 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1060 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1073 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1096 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1112 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1209 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1221 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1306 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1364 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1372 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1445 ();
 sky130_fd_sc_hd__fill_8 FILLER_115_1477 ();
 sky130_fd_sc_hd__fill_4 FILLER_115_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1489 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_81 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_840 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_996 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1032 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1071 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1209 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_116_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1315 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1328 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1332 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1353 ();
 sky130_fd_sc_hd__fill_4 FILLER_116_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1433 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1458 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1460 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1474 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_259 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_861 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_915 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1050 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1105 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1150 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1301 ();
 sky130_fd_sc_hd__fill_4 FILLER_117_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1330 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1346 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_117_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1449 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_297 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_344 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_455 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_488 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_771 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_814 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1068 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1253 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1332 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1355 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1360 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1364 ();
 sky130_fd_sc_hd__fill_4 FILLER_118_1399 ();
 sky130_fd_sc_hd__fill_8 FILLER_118_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1419 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_199 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_207 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_330 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_584 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1086 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1120 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1138 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1207 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1234 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1250 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1267 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1354 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1362 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1378 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1422 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1427 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1435 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_119_1441 ();
 sky130_fd_sc_hd__fill_4 FILLER_119_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_594 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_640 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_652 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_964 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_980 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1013 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1060 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1143 ();
 sky130_fd_sc_hd__fill_4 FILLER_120_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1155 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1298 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1328 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1348 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_120_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1400 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1402 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_320 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1054 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1105 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1151 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1163 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1223 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1344 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1352 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1360 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1368 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1376 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1405 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1425 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1429 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1436 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_121_1469 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1477 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1486 ();
 sky130_fd_sc_hd__fill_4 FILLER_121_1491 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_91 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_105 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_411 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_666 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_682 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_720 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1004 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1072 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1080 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1096 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1184 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1308 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1425 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1432 ();
 sky130_fd_sc_hd__fill_4 FILLER_122_1440 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1444 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1477 ();
 sky130_fd_sc_hd__fill_8 FILLER_122_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1493 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_274 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_532 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_574 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_608 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_693 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_921 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_983 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1072 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1099 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1116 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1124 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1132 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1215 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1219 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1357 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1365 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_123_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_123_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1439 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1496 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_159 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_550 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1074 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1082 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1150 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1169 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1176 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1205 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1213 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1226 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1328 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1357 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1371 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1387 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1395 ();
 sky130_fd_sc_hd__fill_4 FILLER_124_1403 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_124_1448 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1456 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_456 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_545 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1113 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1245 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1282 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1284 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1316 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1336 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1361 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1365 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1388 ();
 sky130_fd_sc_hd__fill_8 FILLER_125_1396 ();
 sky130_fd_sc_hd__fill_4 FILLER_125_1434 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1438 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_130 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_186 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_216 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_224 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_232 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_785 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_817 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_949 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1216 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1226 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1247 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1282 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_126_1297 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1329 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1438 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1450 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1456 ();
 sky130_fd_sc_hd__fill_4 FILLER_126_1465 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_157 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_330 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_464 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_472 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_561 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_638 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_812 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_998 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1006 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1113 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1174 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1342 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1395 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1425 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1433 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1439 ();
 sky130_fd_sc_hd__fill_4 FILLER_127_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1445 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1447 ();
 sky130_fd_sc_hd__fill_8 FILLER_127_1479 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1487 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1489 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_180 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_313 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_604 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1143 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1151 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1161 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1175 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1215 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1256 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1268 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1300 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1314 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1322 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1330 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1338 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1346 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1359 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1370 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1387 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1393 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1432 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1440 ();
 sky130_fd_sc_hd__fill_4 FILLER_128_1448 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1452 ();
 sky130_fd_sc_hd__fill_8 FILLER_128_1460 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1468 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_231 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_390 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_818 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_830 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1121 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1143 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1213 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1285 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1292 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1300 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1308 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1370 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1385 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1396 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1410 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1423 ();
 sky130_fd_sc_hd__fill_8 FILLER_129_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1439 ();
 sky130_fd_sc_hd__fill_4 FILLER_129_1489 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_217 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_262 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_318 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_459 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_467 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_906 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_914 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1249 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1346 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1403 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1409 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_130_1424 ();
 sky130_fd_sc_hd__fill_4 FILLER_130_1464 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1468 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_222 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_452 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_666 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_709 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_752 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1099 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1156 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1225 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1285 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1344 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1346 ();
 sky130_fd_sc_hd__fill_4 FILLER_131_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1407 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_131_1464 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1472 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1474 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_234 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_248 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_322 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_664 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_672 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_835 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1135 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1206 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1222 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1255 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1263 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1298 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1302 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1343 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1360 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1362 ();
 sky130_fd_sc_hd__fill_8 FILLER_132_1372 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1380 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1384 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1386 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_132_1422 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1426 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1428 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1466 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_260 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_576 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_627 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_644 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_709 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1099 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1185 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1209 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1310 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1332 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1376 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1394 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1396 ();
 sky130_fd_sc_hd__fill_8 FILLER_133_1404 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1412 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1436 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1444 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1448 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1452 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1478 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1480 ();
 sky130_fd_sc_hd__fill_4 FILLER_133_1484 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1488 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_334 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_404 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_414 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_595 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_622 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_723 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1113 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1202 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1262 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1356 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1364 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1372 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1380 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1388 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1396 ();
 sky130_fd_sc_hd__fill_4 FILLER_134_1404 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1408 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_134_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1444 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_283 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_616 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_732 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_758 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_870 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_878 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_983 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1118 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1240 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1258 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1267 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1275 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1361 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1385 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1395 ();
 sky130_fd_sc_hd__fill_4 FILLER_135_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1422 ();
 sky130_fd_sc_hd__fill_8 FILLER_135_1432 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1492 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_417 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_633 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_720 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1148 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1253 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1313 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1325 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_136_1427 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1431 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1447 ();
 sky130_fd_sc_hd__fill_8 FILLER_136_1462 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1474 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_312 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_436 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_444 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_507 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_863 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1053 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1065 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1161 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1198 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1357 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1365 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_137_1430 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1438 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1445 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1465 ();
 sky130_fd_sc_hd__fill_4 FILLER_137_1470 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1474 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_174 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_417 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_556 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_654 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_833 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_889 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1140 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1148 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1188 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1196 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1314 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1316 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1346 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1366 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1374 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1400 ();
 sky130_fd_sc_hd__fill_4 FILLER_138_1406 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_138_1438 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1446 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_772 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_930 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_938 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_987 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1110 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1138 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1172 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1180 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1219 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1259 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1283 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1357 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1365 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_139_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1431 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1438 ();
 sky130_fd_sc_hd__fill_8 FILLER_139_1448 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1456 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_286 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_315 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_352 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_395 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_413 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_577 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_994 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1006 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1128 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1144 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1189 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1338 ();
 sky130_fd_sc_hd__fill_4 FILLER_140_1346 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_140_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1462 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_124 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_132 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_140 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_334 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_572 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1163 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1242 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1283 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1312 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1325 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1354 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1368 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1376 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1427 ();
 sky130_fd_sc_hd__fill_4 FILLER_141_1435 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1439 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_141_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1467 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_125 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_483 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_509 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_554 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_605 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_837 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_914 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_967 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1028 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1099 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1103 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1122 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1134 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1186 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1206 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1260 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1309 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1314 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1322 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1370 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1382 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1384 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1427 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1435 ();
 sky130_fd_sc_hd__fill_4 FILLER_142_1445 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1453 ();
 sky130_fd_sc_hd__fill_8 FILLER_142_1461 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_258 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_320 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_328 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_340 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_450 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_692 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_910 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_981 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1076 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1154 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1174 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1286 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1298 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1332 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1354 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1394 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1425 ();
 sky130_fd_sc_hd__fill_4 FILLER_143_1433 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_143_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1462 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1470 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_215 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_493 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_676 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_698 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_953 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1005 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1033 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1065 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1073 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1122 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1197 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1206 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1226 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1237 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1296 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1310 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1324 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1332 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1363 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_144_1430 ();
 sky130_fd_sc_hd__fill_4 FILLER_144_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1446 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1448 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_150 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_946 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_984 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1182 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1190 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1288 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1308 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1316 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1325 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1353 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1399 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1407 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1423 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_145_1454 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1462 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1470 ();
 sky130_fd_sc_hd__fill_4 FILLER_145_1477 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1487 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1489 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_125 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_230 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_326 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_513 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_540 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_862 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_980 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1202 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1210 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1226 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1243 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1245 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1253 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1273 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1323 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1331 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1346 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1372 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1390 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1398 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1402 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1427 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1438 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1442 ();
 sky130_fd_sc_hd__fill_8 FILLER_146_1447 ();
 sky130_fd_sc_hd__fill_4 FILLER_146_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1468 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1474 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_163 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_259 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_286 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_576 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_690 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_865 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1239 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1300 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1302 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1404 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1412 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1420 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1428 ();
 sky130_fd_sc_hd__fill_4 FILLER_147_1436 ();
 sky130_fd_sc_hd__fill_8 FILLER_147_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1461 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_142 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_253 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_394 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_408 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_537 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_597 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_668 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_775 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_787 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1062 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1189 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1206 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1255 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1267 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1272 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1300 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1328 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1336 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1386 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_1394 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1398 ();
 sky130_fd_sc_hd__fill_8 FILLER_148_1402 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1419 ();
 sky130_fd_sc_hd__fill_4 FILLER_148_1448 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1452 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1460 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1468 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_199 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_582 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_621 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_673 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_787 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_867 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_910 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_976 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1099 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1107 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1165 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1230 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_149_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1422 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1430 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1438 ();
 sky130_fd_sc_hd__fill_8 FILLER_149_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1468 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_300 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_403 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_471 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_536 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_592 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_614 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_703 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_707 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1207 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1219 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1246 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1254 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1262 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1266 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1281 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1295 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1334 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1392 ();
 sky130_fd_sc_hd__fill_4 FILLER_150_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_150_1453 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1461 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_401 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_495 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_681 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_718 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_727 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_981 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1146 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1170 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1236 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1248 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1297 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1327 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1352 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1357 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1378 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1398 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1403 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1407 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1420 ();
 sky130_fd_sc_hd__fill_4 FILLER_151_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1433 ();
 sky130_fd_sc_hd__fill_8 FILLER_151_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_477 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_612 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_695 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_710 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1042 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1087 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1104 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1125 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1311 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1320 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1336 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1368 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1376 ();
 sky130_fd_sc_hd__fill_8 FILLER_152_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1408 ();
 sky130_fd_sc_hd__fill_4 FILLER_152_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1415 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1444 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1466 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_325 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_463 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_625 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_754 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_925 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_933 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_979 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_987 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1065 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1216 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1279 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1287 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1295 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1338 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1401 ();
 sky130_fd_sc_hd__fill_8 FILLER_153_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1419 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1430 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1432 ();
 sky130_fd_sc_hd__fill_4 FILLER_153_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_182 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_220 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_240 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_649 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_663 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_966 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1039 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1123 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1204 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1212 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1348 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1355 ();
 sky130_fd_sc_hd__fill_4 FILLER_154_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1369 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1386 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1394 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1413 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1423 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1429 ();
 sky130_fd_sc_hd__fill_8 FILLER_154_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1445 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1474 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_245 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_692 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_724 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_756 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1026 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1038 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1056 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1072 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1117 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1124 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1236 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1293 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1305 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1343 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_155_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1404 ();
 sky130_fd_sc_hd__fill_4 FILLER_155_1417 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1428 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1430 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1438 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_174 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_186 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_242 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_295 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_470 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_495 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_916 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_956 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1022 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1030 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1058 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1076 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1299 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1313 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1369 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1386 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1402 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1409 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1425 ();
 sky130_fd_sc_hd__fill_8 FILLER_156_1433 ();
 sky130_fd_sc_hd__fill_4 FILLER_156_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1445 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1495 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_143 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_353 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_442 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_470 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_716 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_766 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_810 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_814 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_967 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_992 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1041 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1050 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1076 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1095 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1116 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1124 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1154 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1281 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1305 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1336 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1405 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1409 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1414 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1418 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1430 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1432 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_157_1449 ();
 sky130_fd_sc_hd__fill_4 FILLER_157_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1461 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_136 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_360 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_482 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_616 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_770 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_919 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_977 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1088 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1143 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1168 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1188 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1234 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1238 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1315 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1323 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1369 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1377 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1393 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1427 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_158_1460 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1468 ();
 sky130_fd_sc_hd__fill_4 FILLER_158_1471 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1475 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1477 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1484 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1486 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_116 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_336 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_466 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1035 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1039 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1047 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1110 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1170 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1191 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1211 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1237 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1285 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1305 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1310 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1333 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1346 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1354 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1362 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_159_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1399 ();
 sky130_fd_sc_hd__fill_4 FILLER_159_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_135 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_292 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_473 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_682 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_843 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1009 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1026 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1071 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1144 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1158 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1268 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1318 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1328 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1386 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1402 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1420 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1430 ();
 sky130_fd_sc_hd__fill_4 FILLER_160_1438 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1442 ();
 sky130_fd_sc_hd__fill_8 FILLER_160_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1471 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_11 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_36 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_44 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_52 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_214 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_246 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_327 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_487 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_832 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_890 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_980 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1086 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1094 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1208 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1226 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_161_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1394 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1402 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1410 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1412 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_161_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_169 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_184 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_237 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_615 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_769 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_970 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1133 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1303 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1362 ();
 sky130_fd_sc_hd__fill_8 FILLER_162_1370 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1382 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1404 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1408 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1420 ();
 sky130_fd_sc_hd__fill_4 FILLER_162_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1445 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_330 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_338 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_416 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_807 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_919 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_955 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1066 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1251 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1281 ();
 sky130_fd_sc_hd__fill_4 FILLER_163_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_163_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1439 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1455 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1490 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1494 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_304 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_351 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_484 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_515 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_795 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_829 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1010 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1018 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1115 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1178 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1258 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1266 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1270 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1332 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1370 ();
 sky130_fd_sc_hd__fill_8 FILLER_164_1387 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1409 ();
 sky130_fd_sc_hd__fill_4 FILLER_164_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1463 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1468 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1491 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_208 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_257 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_587 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_647 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_728 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_807 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_955 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1025 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1072 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1105 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1117 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1267 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1311 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1342 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1350 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_165_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_165_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1449 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1491 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1496 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_148 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_297 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_319 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_432 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_720 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_796 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_835 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1080 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1206 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1281 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1295 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1374 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1382 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1390 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1398 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1406 ();
 sky130_fd_sc_hd__fill_4 FILLER_166_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_166_1462 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_207 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_238 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_382 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_390 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_454 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_462 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_510 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_570 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_887 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_919 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1123 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1181 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1189 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1282 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1290 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1308 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1335 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1405 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1433 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1439 ();
 sky130_fd_sc_hd__fill_4 FILLER_167_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1466 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1470 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1478 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1482 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1484 ();
 sky130_fd_sc_hd__fill_8 FILLER_167_1488 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_5 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_17 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_593 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_612 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_670 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_735 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_742 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1020 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1089 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1146 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1179 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1205 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1246 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1263 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1289 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1315 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1400 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1408 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1415 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1417 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1433 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1458 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1466 ();
 sky130_fd_sc_hd__fill_8 FILLER_168_1471 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1479 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1483 ();
 sky130_fd_sc_hd__fill_4 FILLER_168_1488 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1492 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_127 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_392 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_465 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_501 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_623 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_653 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_898 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1054 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1167 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1249 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1285 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1387 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1395 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1403 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1427 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1435 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_169_1473 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1481 ();
 sky130_fd_sc_hd__fill_4 FILLER_169_1488 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1492 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_202 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_345 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_720 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_794 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_966 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1057 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1063 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1131 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1161 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1219 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1249 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1301 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1328 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1332 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1382 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1388 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1396 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1400 ();
 sky130_fd_sc_hd__fill_4 FILLER_170_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1440 ();
 sky130_fd_sc_hd__fill_8 FILLER_170_1448 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1469 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_170 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_381 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_430 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_505 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_573 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_675 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_850 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_896 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1030 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1063 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1281 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1333 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1405 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1441 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1474 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1478 ();
 sky130_fd_sc_hd__fill_8 FILLER_171_1482 ();
 sky130_fd_sc_hd__fill_4 FILLER_171_1490 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1494 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_114 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_521 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_594 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_710 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1048 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1270 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1276 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1305 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1327 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1335 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1339 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1416 ();
 sky130_fd_sc_hd__fill_8 FILLER_172_1424 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1432 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1436 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1458 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1460 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1468 ();
 sky130_fd_sc_hd__fill_4 FILLER_172_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_109 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_229 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_274 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_324 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_424 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_440 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_532 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_567 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_581 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_611 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_642 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_844 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_856 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_883 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1170 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1347 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1368 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1376 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_173_1469 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1490 ();
 sky130_fd_sc_hd__fill_4 FILLER_173_1494 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_111 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_166 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_195 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_254 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_262 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_306 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_497 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_521 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_550 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_724 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_928 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_988 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1146 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1189 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1210 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1270 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1272 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1316 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1392 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_174_1479 ();
 sky130_fd_sc_hd__fill_4 FILLER_174_1487 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1491 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_193 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_245 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_283 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_342 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_397 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_567 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_645 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_776 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_872 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1233 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1303 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1326 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1364 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1398 ();
 sky130_fd_sc_hd__fill_8 FILLER_175_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1441 ();
 sky130_fd_sc_hd__fill_4 FILLER_175_1490 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1494 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_115 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_349 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_548 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_662 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_715 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_833 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_978 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1077 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1090 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1130 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1200 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1229 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1242 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1253 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1338 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1383 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1418 ();
 sky130_fd_sc_hd__fill_8 FILLER_176_1471 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1481 ();
 sky130_fd_sc_hd__fill_4 FILLER_176_1494 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1498 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_4 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_18 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_26 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_34 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_42 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_358 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_385 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_483 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_500 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_643 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_694 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_756 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1153 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1180 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1218 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1224 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1232 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1305 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1372 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1407 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1428 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1433 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1439 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1441 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1445 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1471 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1483 ();
 sky130_fd_sc_hd__fill_8 FILLER_177_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_177_1495 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_99 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_171 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_183 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_310 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_717 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_854 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_862 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_910 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1015 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1048 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1055 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1070 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1119 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1158 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1180 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1188 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1206 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1246 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1281 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1297 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1309 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1382 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1466 ();
 sky130_fd_sc_hd__fill_8 FILLER_178_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1482 ();
 sky130_fd_sc_hd__fill_4 FILLER_178_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1496 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_113 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_452 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_539 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_550 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_619 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_712 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_874 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_930 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_952 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1073 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1099 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1198 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1224 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1232 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1240 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1248 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1280 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1300 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1312 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1321 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1396 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1404 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1412 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1455 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1463 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_179_1479 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_179_1492 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_121 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_600 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_637 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_653 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_726 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_862 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1015 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1066 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1074 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1197 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1253 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1279 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1305 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1313 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1377 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1390 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1437 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1478 ();
 sky130_fd_sc_hd__fill_8 FILLER_180_1486 ();
 sky130_fd_sc_hd__fill_4 FILLER_180_1494 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_168 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_176 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_560 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_620 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_628 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_934 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1066 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1143 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1180 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1285 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1305 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1316 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1346 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1354 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1381 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1389 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1393 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1400 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1410 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1414 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1439 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1445 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1452 ();
 sky130_fd_sc_hd__fill_8 FILLER_181_1480 ();
 sky130_fd_sc_hd__fill_4 FILLER_181_1488 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_109 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_377 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_633 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_835 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_847 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_989 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1072 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1180 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1218 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1226 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1231 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1243 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1278 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1286 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1355 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1360 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1362 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1379 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1387 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1391 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1396 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1444 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1453 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1461 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1471 ();
 sky130_fd_sc_hd__fill_4 FILLER_182_1479 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1483 ();
 sky130_fd_sc_hd__fill_8 FILLER_182_1488 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_93 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_112 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_178 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_356 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_433 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_452 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_572 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_743 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_786 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_863 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_915 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_934 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_985 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1039 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1102 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1189 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1209 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1264 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1272 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1280 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1319 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1321 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1327 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1342 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1344 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1354 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1362 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1459 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1467 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1475 ();
 sky130_fd_sc_hd__fill_8 FILLER_183_1483 ();
 sky130_fd_sc_hd__fill_4 FILLER_183_1491 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_196 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_292 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_573 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_663 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_714 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_730 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1017 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1102 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1142 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1237 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1249 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1376 ();
 sky130_fd_sc_hd__fill_4 FILLER_184_1384 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1388 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1390 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1435 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1445 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1471 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_184_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1491 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_101 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_285 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_293 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_510 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_966 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_992 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1043 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1159 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1176 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1237 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1278 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1304 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1312 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1331 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1339 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1365 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1403 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1408 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1416 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1424 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1438 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1461 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_185_1477 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1485 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1489 ();
 sky130_fd_sc_hd__fill_4 FILLER_185_1494 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1498 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_112 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_120 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_128 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_275 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_587 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_595 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_715 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_735 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_853 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1007 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1030 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1098 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1129 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1162 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1210 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1223 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1238 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1264 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1268 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1270 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1310 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1325 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1341 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1367 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1408 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1418 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1422 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1454 ();
 sky130_fd_sc_hd__fill_8 FILLER_186_1462 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1471 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1475 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1477 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1481 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1485 ();
 sky130_fd_sc_hd__fill_4 FILLER_186_1492 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_276 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_543 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_586 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_637 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_677 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_701 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_948 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1047 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1064 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1072 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1275 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1307 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1324 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1332 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1336 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1346 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1354 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1370 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1389 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1403 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1428 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1432 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1454 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1462 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1470 ();
 sky130_fd_sc_hd__fill_8 FILLER_187_1475 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1487 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1489 ();
 sky130_fd_sc_hd__fill_4 FILLER_187_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_146 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_173 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_350 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_409 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_466 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_487 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_547 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_563 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_655 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_667 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_784 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_792 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_808 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_922 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1130 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1146 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1261 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1273 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1295 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1338 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1346 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1382 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1386 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1388 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1392 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1400 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1402 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1465 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1471 ();
 sky130_fd_sc_hd__fill_4 FILLER_188_1479 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1483 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1485 ();
 sky130_fd_sc_hd__fill_8 FILLER_188_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1497 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_7 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_15 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_23 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_154 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_212 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_230 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_336 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_387 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_549 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_565 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_609 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_665 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_737 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1085 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1101 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1145 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1188 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1216 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1234 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1242 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1271 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1306 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1318 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1344 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1352 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1356 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_189_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1457 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1482 ();
 sky130_fd_sc_hd__fill_4 FILLER_189_1489 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1493 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_285 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_546 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_620 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_647 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_791 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_868 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1124 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1221 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1228 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1260 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1268 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1289 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1298 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1310 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_190_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1349 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1353 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1362 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1364 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1372 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1380 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1382 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1427 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1435 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1443 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1445 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1475 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1483 ();
 sky130_fd_sc_hd__fill_8 FILLER_190_1491 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_4 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_17 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_25 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_119 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_206 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_298 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_326 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_559 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_584 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_641 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_679 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_687 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_695 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_913 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1249 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1253 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1265 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1283 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1287 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1305 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1366 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1392 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1400 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1408 ();
 sky130_fd_sc_hd__fill_4 FILLER_191_1419 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1425 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_191_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1497 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_0 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_123 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_138 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_146 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_221 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_308 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_441 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_529 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_537 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_821 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_939 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1039 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1046 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1146 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1155 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1295 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1351 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1423 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1431 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_192_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_192_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_33 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_41 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_341 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_648 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1040 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1063 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1126 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1132 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1209 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1253 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1261 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1265 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1316 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1342 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1350 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1362 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1401 ();
 sky130_fd_sc_hd__fill_4 FILLER_193_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_193_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_498 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_506 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_629 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_639 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_851 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1075 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1149 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1166 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1186 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1194 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1210 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1267 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1294 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1305 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1323 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1395 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1411 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1450 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1458 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1466 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_194_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_194_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_214 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_313 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_321 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_337 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_345 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_464 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_547 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_578 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_643 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_667 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_671 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_867 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_947 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_973 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1006 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1057 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1078 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1117 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1172 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1196 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1224 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1269 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1278 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1280 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1301 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1323 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1351 ();
 sky130_fd_sc_hd__fill_4 FILLER_195_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1378 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1385 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1393 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1409 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1411 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_195_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_290 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_343 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_407 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_453 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_496 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_540 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_634 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_829 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_837 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1004 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1092 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1115 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1133 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1177 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1211 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1238 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1279 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1338 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_1344 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1348 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1360 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1372 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1394 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1402 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1432 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1440 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1448 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1456 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_1464 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1468 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_196_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_196_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_3 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_11 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_19 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_129 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_141 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_228 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_232 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_318 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_346 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_443 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_468 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_499 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_623 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_656 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_745 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_761 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_896 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_941 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1068 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1083 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1141 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1155 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1176 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1227 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1266 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1273 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1300 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1313 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1366 ();
 sky130_fd_sc_hd__fill_4 FILLER_197_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1378 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1432 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_197_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_139 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_282 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_294 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_353 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_597 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_613 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_655 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1125 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1158 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1166 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1193 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1197 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1205 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1242 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1250 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1299 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1316 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1339 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1349 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1363 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1395 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1403 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_198_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_198_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_134 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_359 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_382 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_507 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_535 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_565 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_581 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_763 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_935 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_987 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1039 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_1100 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1112 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1123 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1185 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1209 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1288 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1366 ();
 sky130_fd_sc_hd__fill_4 FILLER_199_1374 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1378 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1405 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_199_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_373 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_531 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_610 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_651 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_815 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_858 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_866 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_986 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_999 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1084 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1145 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1267 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1291 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1303 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1332 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1340 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1348 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1408 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_200_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_200_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_176 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_193 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_213 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_319 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_516 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_524 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_785 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1073 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1100 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1174 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1201 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1213 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1220 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1232 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1240 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1287 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_1295 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1343 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_201_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1379 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1407 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1415 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1423 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_201_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_131 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_357 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_403 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_430 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_475 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_686 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_717 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1039 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1057 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1074 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1121 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1129 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1186 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1198 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1206 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1259 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1280 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1291 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1329 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1346 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1358 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1366 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1374 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1382 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1390 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1398 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1406 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_202_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_202_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_278 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_373 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_453 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_503 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_576 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_683 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_702 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_726 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_731 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_739 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_797 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_974 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_996 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1039 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1112 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1230 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1245 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_1253 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_203_1277 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1319 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1339 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1347 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1355 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1363 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_203_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_219 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_289 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_636 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_786 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_794 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_817 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_913 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_960 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1026 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1060 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1074 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1108 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1123 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1136 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1146 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1214 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1234 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1248 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1264 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1272 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1276 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1278 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1286 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1291 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1295 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1302 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1310 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1321 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1325 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1342 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_204_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_204_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_236 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_253 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_273 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_445 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_528 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_556 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_598 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_915 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1021 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1039 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1047 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1090 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1098 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1106 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1114 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1122 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1138 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1248 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1269 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1297 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1305 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1328 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1336 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1344 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1352 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1360 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1368 ();
 sky130_fd_sc_hd__fill_4 FILLER_205_1376 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_205_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_10 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_139 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_191 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_233 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_388 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_411 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_427 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_611 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_759 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_865 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_913 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_965 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1073 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1154 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_1162 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1182 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1200 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1258 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1266 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1274 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1282 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_206_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_206_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_8 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_27 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_35 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_43 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_154 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_307 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_311 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_323 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_439 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_599 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_789 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_919 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1010 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1123 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1138 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1156 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_207_1243 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_207_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1497 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_0 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_9 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_215 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_479 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_552 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_557 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_569 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_605 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_679 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_802 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_903 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_918 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1014 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1022 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1038 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1069 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1130 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1184 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1192 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1200 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1248 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1256 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1264 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1272 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1280 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1288 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_208_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_208_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_20 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_204 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_330 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_437 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_517 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_585 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_825 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_880 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_888 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_994 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1059 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1071 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1085 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1094 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1108 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_1116 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1125 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1174 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1199 ();
 sky130_fd_sc_hd__fill_4 FILLER_209_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1207 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1239 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_209_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_160 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_172 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_217 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_248 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_436 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_462 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_602 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_895 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_931 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1111 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1173 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_1179 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1237 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1257 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_210_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_210_1495 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_228 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_236 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_358 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_524 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_593 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_632 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1008 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_1016 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1041 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1049 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1110 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1139 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_211_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_211_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1497 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_2 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_13 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_29 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_155 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_172 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_198 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_206 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_233 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_449 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_460 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_488 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_517 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_711 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_733 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_767 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_928 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1051 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1070 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1084 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1160 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1228 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1235 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_212_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_212_1495 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_0 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_2 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_6 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_14 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_22 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_30 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_38 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_46 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_58 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_225 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_309 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_356 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_425 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_497 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_567 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_698 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_729 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_793 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_919 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1092 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1106 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1152 ();
 sky130_fd_sc_hd__fill_4 FILLER_213_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1178 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1246 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1251 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_213_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_149 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_157 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_289 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_317 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_429 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_437 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_544 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_566 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_575 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_594 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_602 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_732 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_736 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_805 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1020 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1025 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1033 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1077 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1109 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_214_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_214_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_155 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_188 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_404 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_467 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_505 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_609 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_646 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_688 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_810 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_848 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_938 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1027 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1050 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1062 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1079 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1093 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1144 ();
 sky130_fd_sc_hd__fill_4 FILLER_215_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_215_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_208 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_211 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_226 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_402 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_414 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_546 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_589 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_613 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_643 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_662 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_753 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_888 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_900 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_980 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_986 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1019 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1088 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1147 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1185 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1249 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1257 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1265 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1273 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_216_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_216_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_299 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_330 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_569 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_617 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_826 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_849 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_890 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_901 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_915 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_979 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1029 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1050 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1083 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1110 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1134 ();
 sky130_fd_sc_hd__fill_4 FILLER_217_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1183 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1236 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1244 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1252 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_217_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_237 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_260 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_363 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_424 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_508 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_515 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_527 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_555 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_664 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_774 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_801 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_819 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_915 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1003 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1020 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1028 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_1036 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1128 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1147 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1171 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_1178 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1214 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1222 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_218_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_218_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_223 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_263 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_396 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_412 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_425 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_584 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_700 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_752 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_772 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_936 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1005 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1087 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_1095 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1117 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1129 ();
 sky130_fd_sc_hd__fill_4 FILLER_219_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_219_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_269 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_378 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_391 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_446 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_529 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_543 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_610 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_734 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_742 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_775 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_907 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_923 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1033 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1075 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1140 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1148 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1156 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1168 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_220_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_220_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_189 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_203 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_322 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_369 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_429 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_441 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_461 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_472 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_625 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_641 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_729 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_755 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_807 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_838 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_965 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_970 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_978 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1081 ();
 sky130_fd_sc_hd__fill_4 FILLER_221_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1132 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_221_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_161 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_190 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_316 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_389 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_534 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_568 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_615 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_877 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_943 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1009 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1130 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1138 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1146 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1154 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1162 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_222_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_222_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_165 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_178 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_323 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_396 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_489 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_658 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_697 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_725 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_730 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_738 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_750 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_799 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_859 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_867 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_884 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_892 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_922 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_934 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_979 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1004 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1012 ();
 sky130_fd_sc_hd__fill_4 FILLER_223_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_223_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_151 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_190 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_250 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_266 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_335 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_438 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_446 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_457 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_465 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_591 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_650 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_699 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_707 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_771 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_790 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_802 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1016 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1024 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1032 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_224_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_224_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_247 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_255 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_365 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_380 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_416 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_421 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_455 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_548 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_559 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_658 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_750 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_806 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_845 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_891 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_969 ();
 sky130_fd_sc_hd__fill_4 FILLER_225_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_225_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_239 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_268 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_349 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_431 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_676 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_697 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_701 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_709 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_727 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_746 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_769 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_816 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_824 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_832 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_875 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_226_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_226_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_145 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_333 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_478 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_485 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_549 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_558 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_806 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_937 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_945 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_959 ();
 sky130_fd_sc_hd__fill_4 FILLER_227_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_227_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_287 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_355 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_367 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_456 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_469 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_494 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_502 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_589 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_677 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_748 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_809 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_842 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_862 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_929 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_991 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1037 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_228_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_228_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_153 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_165 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_205 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_244 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_307 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_342 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_439 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_501 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_513 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_627 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_652 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_716 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_725 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_779 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_787 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_806 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_818 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_822 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_838 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_863 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_952 ();
 sky130_fd_sc_hd__fill_4 FILLER_229_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_229_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_169 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_194 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_202 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_293 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_305 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_367 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_449 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_475 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_523 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_554 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_562 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_578 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_639 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_782 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_834 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_897 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_968 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_230_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_230_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_179 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_185 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_379 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_447 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_526 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_553 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_669 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_940 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_948 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_956 ();
 sky130_fd_sc_hd__fill_4 FILLER_231_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_231_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_229 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_258 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_266 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_294 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_306 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_331 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_343 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_381 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_398 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_579 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_693 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_753 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_837 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_875 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_953 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1027 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1035 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_232_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_232_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_222 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_296 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_347 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_404 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_412 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_454 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_458 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_526 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_545 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_564 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_820 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_836 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_952 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_979 ();
 sky130_fd_sc_hd__fill_4 FILLER_233_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_233_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_185 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_370 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_427 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_480 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_519 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_631 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_675 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_689 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_691 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_731 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_757 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_761 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_777 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_853 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_926 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1020 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_234_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_234_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_238 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_247 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_281 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_348 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_405 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_419 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_476 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_481 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_544 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_564 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_572 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_580 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_684 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_704 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_712 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_737 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_859 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_895 ();
 sky130_fd_sc_hd__fill_4 FILLER_235_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_997 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_235_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_175 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_187 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_223 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_277 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_339 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_431 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_568 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_571 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_640 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_648 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_686 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_722 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_749 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_770 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_782 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_905 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_958 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_970 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1012 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1020 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1028 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1036 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1048 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_236_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_236_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_181 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_265 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_379 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_460 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_489 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_527 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_539 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_603 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_705 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_721 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_741 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_755 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_839 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_907 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_237_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_237_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_209 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_279 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_302 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_409 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_435 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_477 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_491 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_519 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_628 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_635 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_730 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_783 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_889 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_897 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_911 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_955 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_988 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_238_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_238_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_271 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_303 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_415 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_479 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_491 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_514 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_557 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_619 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_659 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_661 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_673 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_765 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_861 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_909 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_961 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_973 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_990 ();
 sky130_fd_sc_hd__fill_4 FILLER_239_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1002 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1018 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_239_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_235 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_264 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_408 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_428 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_536 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_562 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_571 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_583 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_626 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_689 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_703 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_746 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_783 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_837 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_871 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_883 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_975 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_240_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_240_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_251 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_310 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_365 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_418 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_445 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_478 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_481 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_511 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_525 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_541 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_585 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_599 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_607 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_634 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_685 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_705 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_841 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_868 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_927 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_935 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_943 ();
 sky130_fd_sc_hd__fill_4 FILLER_241_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_967 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_241_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_242_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_243 ();
 sky130_fd_sc_hd__fill_4 FILLER_242_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_255 ();
 sky130_fd_sc_hd__fill_4 FILLER_242_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_268 ();
 sky130_fd_sc_hd__fill_4 FILLER_242_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_275 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_338 ();
 sky130_fd_sc_hd__fill_4 FILLER_242_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_451 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_551 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_592 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_629 ();
 sky130_fd_sc_hd__fill_4 FILLER_242_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_671 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_757 ();
 sky130_fd_sc_hd__fill_4 FILLER_242_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_791 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_811 ();
 sky130_fd_sc_hd__fill_4 FILLER_242_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_823 ();
 sky130_fd_sc_hd__fill_4 FILLER_242_866 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_242_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_242_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_243_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_282 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_298 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_301 ();
 sky130_fd_sc_hd__fill_4 FILLER_243_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_394 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_448 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_538 ();
 sky130_fd_sc_hd__fill_4 FILLER_243_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_583 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_588 ();
 sky130_fd_sc_hd__fill_4 FILLER_243_596 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_706 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_719 ();
 sky130_fd_sc_hd__fill_4 FILLER_243_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_243_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_800 ();
 sky130_fd_sc_hd__fill_4 FILLER_243_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_823 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_828 ();
 sky130_fd_sc_hd__fill_4 FILLER_243_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_885 ();
 sky130_fd_sc_hd__fill_4 FILLER_243_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_899 ();
 sky130_fd_sc_hd__fill_4 FILLER_243_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_910 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_918 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_926 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_934 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_942 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_958 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_243_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_244_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_314 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_388 ();
 sky130_fd_sc_hd__fill_4 FILLER_244_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_448 ();
 sky130_fd_sc_hd__fill_4 FILLER_244_451 ();
 sky130_fd_sc_hd__fill_4 FILLER_244_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_508 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_244_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_523 ();
 sky130_fd_sc_hd__fill_4 FILLER_244_566 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_579 ();
 sky130_fd_sc_hd__fill_4 FILLER_244_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_636 ();
 sky130_fd_sc_hd__fill_4 FILLER_244_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_749 ();
 sky130_fd_sc_hd__fill_4 FILLER_244_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_879 ();
 sky130_fd_sc_hd__fill_4 FILLER_244_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_891 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_905 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_244_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_244_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_244_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_245_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_245_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_460 ();
 sky130_fd_sc_hd__fill_4 FILLER_245_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_485 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_541 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_586 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_598 ();
 sky130_fd_sc_hd__fill_4 FILLER_245_601 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_659 ();
 sky130_fd_sc_hd__fill_4 FILLER_245_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_665 ();
 sky130_fd_sc_hd__fill_4 FILLER_245_708 ();
 sky130_fd_sc_hd__fill_4 FILLER_245_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_778 ();
 sky130_fd_sc_hd__fill_4 FILLER_245_788 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_795 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_803 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_827 ();
 sky130_fd_sc_hd__fill_4 FILLER_245_836 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_245_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_246_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_329 ();
 sky130_fd_sc_hd__fill_4 FILLER_246_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_335 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_246_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_375 ();
 sky130_fd_sc_hd__fill_4 FILLER_246_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_423 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_442 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_518 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_603 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_631 ();
 sky130_fd_sc_hd__fill_4 FILLER_246_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_688 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_748 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_751 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_759 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_798 ();
 sky130_fd_sc_hd__fill_4 FILLER_246_806 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_855 ();
 sky130_fd_sc_hd__fill_4 FILLER_246_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_877 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_885 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_893 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_246_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_246_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_246_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_247_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_395 ();
 sky130_fd_sc_hd__fill_4 FILLER_247_421 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_443 ();
 sky130_fd_sc_hd__fill_4 FILLER_247_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_538 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_651 ();
 sky130_fd_sc_hd__fill_4 FILLER_247_656 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_767 ();
 sky130_fd_sc_hd__fill_4 FILLER_247_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_779 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_247_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_248_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_399 ();
 sky130_fd_sc_hd__fill_4 FILLER_248_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_415 ();
 sky130_fd_sc_hd__fill_4 FILLER_248_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_459 ();
 sky130_fd_sc_hd__fill_4 FILLER_248_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_509 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_511 ();
 sky130_fd_sc_hd__fill_4 FILLER_248_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_551 ();
 sky130_fd_sc_hd__fill_4 FILLER_248_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_575 ();
 sky130_fd_sc_hd__fill_4 FILLER_248_622 ();
 sky130_fd_sc_hd__fill_4 FILLER_248_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_635 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_691 ();
 sky130_fd_sc_hd__fill_4 FILLER_248_699 ();
 sky130_fd_sc_hd__fill_4 FILLER_248_706 ();
 sky130_fd_sc_hd__fill_4 FILLER_248_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_717 ();
 sky130_fd_sc_hd__fill_4 FILLER_248_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_758 ();
 sky130_fd_sc_hd__fill_4 FILLER_248_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_799 ();
 sky130_fd_sc_hd__fill_4 FILLER_248_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_989 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1067 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1075 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1083 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1091 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_248_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_248_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_249_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_241 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_257 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_265 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_273 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_281 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_377 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_385 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_393 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_401 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_419 ();
 sky130_fd_sc_hd__fill_4 FILLER_249_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_492 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_525 ();
 sky130_fd_sc_hd__fill_4 FILLER_249_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_249_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_672 ();
 sky130_fd_sc_hd__fill_4 FILLER_249_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_718 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_762 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_778 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_813 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_821 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_881 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_899 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_917 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_925 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_959 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_961 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_969 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_977 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_985 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_993 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1001 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1019 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1021 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1029 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1037 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1045 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1053 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1061 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_249_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_250_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_47 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_55 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_63 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_71 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_107 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_115 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_123 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_131 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_167 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_175 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_183 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_191 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_227 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_235 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_243 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_251 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_269 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_271 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_279 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_287 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_295 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_303 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_311 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_329 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_331 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_339 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_347 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_355 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_363 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_371 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_389 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_407 ();
 sky130_fd_sc_hd__fill_4 FILLER_250_626 ();
 sky130_fd_sc_hd__fill_4 FILLER_250_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_764 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_793 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_809 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_811 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_819 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_827 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_835 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_843 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_851 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_869 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_871 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_879 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_887 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_895 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_903 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_911 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_931 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_939 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_947 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_955 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_963 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_971 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_982 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_991 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_999 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1007 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1015 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1023 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1031 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1055 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1063 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1071 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1087 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1095 ();
 sky130_fd_sc_hd__fill_4 FILLER_250_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1127 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1135 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1143 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1151 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1187 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1195 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1203 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1211 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1247 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1255 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1263 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1271 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1279 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1307 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1315 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1323 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1331 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1339 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1367 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1375 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1383 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1391 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1427 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1435 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1443 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1451 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_1467 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_250_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_250_1495 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_16 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_24 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_32 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_40 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_48 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_56 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_77 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_85 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_93 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_101 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_137 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_145 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_153 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_161 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_197 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_205 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_213 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_221 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_239 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_241 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_249 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_256 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_264 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_272 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_280 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_288 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_296 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_309 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_317 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_325 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_333 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_341 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_359 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_361 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_369 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_376 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_384 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_391 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_399 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_423 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_601 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_617 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_621 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_661 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_669 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_685 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_719 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_721 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_763 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_775 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_781 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_789 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_797 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_805 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_813 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_825 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_857 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_865 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_873 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_881 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_898 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_901 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_909 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_917 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_929 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_933 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_941 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_968 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_976 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_980 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_987 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_995 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1003 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1039 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1043 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1051 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1059 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1067 ();
 sky130_fd_sc_hd__fill_4 FILLER_251_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1097 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1105 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1113 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1121 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1157 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1165 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1173 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1181 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1217 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1225 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1233 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1241 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1249 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1277 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1285 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1293 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1301 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1309 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1337 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1345 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1353 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1361 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1397 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1405 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1413 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1421 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_1437 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1457 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1465 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1473 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1481 ();
 sky130_fd_sc_hd__fill_8 FILLER_251_1489 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_1497 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_0 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_8 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_16 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_28 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_31 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_39 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_47 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_59 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_61 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_69 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_77 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_89 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_91 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_99 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_107 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_119 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_121 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_129 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_137 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_149 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_151 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_159 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_167 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_179 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_181 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_189 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_197 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_209 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_211 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_219 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_227 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_249 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_291 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_299 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_301 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_312 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_328 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_344 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_352 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_361 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_380 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_649 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_678 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_702 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_751 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_768 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_776 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_781 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_839 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_841 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_849 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_857 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_869 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_886 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_903 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_907 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_923 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_937 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_951 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1049 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1057 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1065 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1079 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1081 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1089 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1097 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1109 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1111 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1119 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1127 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1139 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1141 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1149 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1157 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1169 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1171 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1179 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1187 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1199 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1201 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1209 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1217 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1229 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1231 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1239 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1247 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1259 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1261 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1269 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1277 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1289 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1291 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1299 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1307 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1319 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1321 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1329 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1337 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1349 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1351 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1359 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1367 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1379 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1381 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1389 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1397 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_1405 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1409 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1411 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1419 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1427 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_1435 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1439 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1441 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1449 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1457 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_1465 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1469 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1471 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1479 ();
 sky130_fd_sc_hd__fill_8 FILLER_252_1487 ();
 sky130_fd_sc_hd__fill_4 FILLER_252_1495 ();
endmodule
